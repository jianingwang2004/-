
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/04/08 14:43:44
// Design Name: 
// Module Name: CPU
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
`define    PC_INIT      32'H1c000000
`define    HALT_INST    32'H80000000
module CPU (
    input                   [ 0 : 0]            clk,
    input                   [ 0 : 0]            rst,

    input                   [ 0 : 0]            global_en,

/* ------------------------------ Memory (inst) ----------------------------- */
    output                  [31 : 0]            imem_raddr,
    input                   [31 : 0]            imem_rdata,

/* ------------------------------ Memory (data) ----------------------------- */
    input                   [31 : 0]            dmem_rdata,
    output                  [ 0 : 0]            dmem_we,
    output                  [31 : 0]            dmem_addr,
    output                  [31 : 0]            dmem_wdata,

/* ---------------------------------- Debug --------------------------------- */
    output                  [ 0 : 0]            commit,
    output                  [31 : 0]            commit_pc,
    output                  [31 : 0]            commit_inst,
    output                  [ 0 : 0]            commit_halt,
    output                  [ 0 : 0]            commit_reg_we,
    output                  [ 4 : 0]            commit_reg_wa,
    output                  [31 : 0]            commit_reg_wd,
    output                  [ 0 : 0]            commit_dmem_we,
    output                  [31 : 0]            commit_dmem_wa,
    output                  [31 : 0]            commit_dmem_wd,

    input                   [ 4 : 0]            debug_reg_ra,
    output                  [31 : 0]            debug_reg_rd
);

//for PC/NPC_mux
wire [ 1 : 0]     npc_sel;
wire [31 : 0]      npc_ex;
assign imem_raddr = pc_if;

//for IF/ID
wire [31 : 0]   pcadd4_if;
wire [31 : 0]   pcadd4_id;
wire [31 : 0]       pc_if;	
wire [31 : 0]       pc_id;
wire [31 : 0]     inst_id;
wire [ 0 : 0] 	commit_if;
wire [ 0 : 0]	commit_id;
wire [ 0 : 0]       stall;
wire [ 0 : 0]       flush;
assign	stall 	  =  1'b0;
assign 	commit_if =  1'b1;

PC my_pc (
    .clk    (        clk),
    .rst    (        rst),
    .en     (  global_en),    // �� global_en Ϊ�ߵ�ƽʱ��PC �Ż���£�CPU �Ż�ִ��ָ�
    .npc    (     npc_ex),
    .pc     (      pc_if)
);

ADD4 adder(
    .a      (	   pc_if),
    .b      (      32'd4),
    .c      (  pcadd4_if)
);

Intersegment_REG IF_ID(
    .clk		(            clk),
    .rst		(            rst),
    .en			(      global_en),
    .stall		(          stall),
    .flush		(          flush),
      
    .pcadd4_in		(      pcadd4_if),
    .pcadd4_out		(      pcadd4_id),
    .pc_in		(          pc_if),
    .pc_out		(          pc_id),
    .inst_in		(     imem_rdata),
    .inst_out		(        inst_id),
    .commit_in		(      commit_if),
    .commit_out		(      commit_id),
      
    .imm_in		(	   32'd0),
    .imm_out		(		),
    .rf_wa_in		(           5'd0),
    .rf_wa_out		(		),
    .rf_rd0_in		(          32'd0),
    .rf_rd0_out		(		),
    .rf_rd1_in		(          32'd0),
    .rf_rd1_out		(		),
    .rf_we_in		(           1'd0),
    .rf_we_out		(		),
    .rf_wd_sel_in	(           2'd0),
    .rf_wd_sel_out	(		),
    .alu_op_in		(           5'd0),
    .alu_op_out		(		),
    .alu_src0_sel_in	(           1'd0),
    .alu_src0_sel_out	(		),
    .alu_src1_sel_in	(           1'd0),
    .alu_src1_sel_out	(		),
    .dmem_access_in	(           4'd0),
    .dmem_access_out	(		),
    .br_type_in		(           4'd0),
    .br_type_out	(		),
    
    .alu_res_in		(          32'd0),
    .alu_res_out	(		),
            
    .dmem_rd_out_in	(          32'd0),
    .dmem_rd_out_out	(		),
    .dmem_wdata_in	(          32'd0),
    .dmem_wdata_out	(		),
    .dmem_we_in		(           1'd0),
    .dmem_we_out	(		)
);

//for decoder
wire [ 4 : 0]          rf_ra0_id;
wire [ 4 : 0]          rf_ra1_id;


//for ID/EX
wire [31 : 0]          pcadd4_ex;
wire [31 : 0]              pc_ex;
wire [31 : 0]            inst_ex;
wire [ 0 : 0] 	       commit_ex;
wire [31 : 0]             imm_id;
wire [31 : 0]             imm_ex;
wire [ 4 : 0]           rf_wa_id;
wire [ 4 : 0]           rf_wa_ex;
wire [31 : 0]          rf_rd0_id;
wire [31 : 0]          rf_rd0_ex;
wire [31 : 0]          rf_rd1_id;
wire [31 : 0]          rf_rd1_ex;
wire [ 0 : 0]           rf_we_id;
wire [ 0 : 0]           rf_we_ex;
wire [ 1 : 0]       rf_wd_sel_id;
wire [ 1 : 0]       rf_wd_sel_ex;
wire [ 4 : 0]          alu_op_id;
wire [ 4 : 0]          alu_op_ex;
wire [ 0 : 0]    alu_src0_sel_id;
wire [ 0 : 0]    alu_src0_sel_ex;
wire [ 0 : 0]    alu_src1_sel_id;
wire [ 0 : 0]    alu_src1_sel_ex;
wire [ 3 : 0]     dmem_access_id;
wire [ 3 : 0]     dmem_access_ex;
wire [ 3 : 0]         br_type_id;
wire [ 3 : 0]         br_type_ex;
wire [ 0 : 0]         dmem_we_id;
wire [ 0 : 0]         dmem_we_ex;
wire [31 : 0]           rf_wd_wb;
DECODE decode(
    .inst		(	 inst_id),
    .alu_op		(      alu_op_id),
    .dmem_access	( dmem_access_id),
    .imm		(         imm_id),
    .rf_ra0		(      rf_ra0_id),
    .rf_ra1		(      rf_ra1_id),
    .rf_wa		(	rf_wa_id),
    .rf_we		(	rf_we_id),
    .rf_wd_sel		(   rf_wd_sel_id),
    .alu_src0_sel	(alu_src0_sel_id),
    .alu_src1_sel	(alu_src1_sel_id),
    .br_type		(     br_type_id),
    .dmem_we		(     dmem_we_id)
    );
    
REGFILE regfile(
    .clk		(            clk),
    .rf_ra0		(      rf_ra0_id),
    .rf_ra1		(      rf_ra1_id),
    .dbg_reg_ra		(   debug_reg_ra), 
    .rf_wa		(       rf_wa_wb),
    .rf_we		(       rf_we_wb),
    .rf_wd		(       rf_wd_wb),
    .rf_rd0		(      rf_rd0_id),
    .rf_rd1		(      rf_rd1_id),
    .dbg_reg_rd		(   debug_reg_rd)
);

Intersegment_REG ID_EX(
    .clk		(            clk),
    .rst		(            rst),
    .en			(      global_en),
    .stall		(          stall),
    .flush		(          flush),
      
    .pcadd4_in		(      pcadd4_id),
    .pcadd4_out		(      pcadd4_ex),
    .pc_in		(          pc_id),
    .pc_out		(          pc_ex),
    .inst_in		(        inst_id),
    .inst_out		(        inst_ex),
    .commit_in		(      commit_id),
    .commit_out		(      commit_ex),
      
    .imm_in		(	  imm_id),
    .imm_out		(      	  imm_ex),
    .rf_wa_in		(       rf_wa_id),
    .rf_wa_out		(	rf_wa_ex),
    .rf_rd0_in		(      rf_rd0_id),
    .rf_rd0_out		(      rf_rd0_ex),
    .rf_rd1_in		(      rf_rd1_id),
    .rf_rd1_out		(      rf_rd1_ex),
    .rf_we_in		(       rf_we_id),
    .rf_we_out		(       rf_we_ex),
    .rf_wd_sel_in	(   rf_wd_sel_id),
    .rf_wd_sel_out	(   rf_wd_sel_ex),
    .alu_op_in		(      alu_op_id),
    .alu_op_out		(      alu_op_ex),
    .alu_src0_sel_in	(alu_src0_sel_id),
    .alu_src0_sel_out	(alu_src0_sel_ex),
    .alu_src1_sel_in	(alu_src1_sel_id),
    .alu_src1_sel_out	(alu_src1_sel_ex),
    .dmem_access_in	( dmem_access_id),
    .dmem_access_out	( dmem_access_ex),
    .br_type_in		(     br_type_id),
    .br_type_out	(     br_type_ex),
    
    .alu_res_in		(          32'd0),
    .alu_res_out	(		),
            
    .dmem_rd_out_in	(          32'd0),
    .dmem_rd_out_out	(		),
    .dmem_wdata_in	(          32'd0),
    .dmem_wdata_out	(		),
    .dmem_we_in		(     dmem_we_id),
    .dmem_we_out	(     dmem_we_ex)
);

//for alu
wire [31 : 0]   alu_src0_ex;
wire [31 : 0]   alu_src1_ex;

//for EX/MEM
assign flush = (npc_sel == 2'b01) ? 1'b1 : 1'b0;
wire [31 : 0]          pcadd4_mem;
wire [31 : 0]              pc_mem;
wire [31 : 0]            inst_mem;
wire [ 0 : 0]          commit_mem;
wire [31 : 0]             imm_mem;
wire [ 4 : 0]           rf_wa_mem;
wire [31 : 0]          rf_rd0_mem;
wire [31 : 0]          rf_rd1_mem;
wire [ 0 : 0]           rf_we_mem;
wire [ 1 : 0]       rf_wd_sel_mem;
wire [ 4 : 0]          alu_op_mem;
wire [ 0 : 0]    alu_src0_sel_mem;
wire [ 0 : 0]    alu_src1_sel_mem;
wire [ 3 : 0]     dmem_access_mem;
wire [ 3 : 0]         br_type_mem;
wire [ 0 : 0]         dmem_we_mem;
wire [31 : 0]          alu_res_ex;
wire [31 : 0]         alu_res_mem;


BRANCH branch(
    .br_type	(     br_type_ex),
    .br_src0	(      rf_rd0_ex),
    .br_src1	(      rf_rd1_ex),
    .npc_sel	(        npc_sel)
);

MUX mux0(
    .src0	(      rf_rd0_ex), 
    .src1	(          pc_ex),
    .sel	(alu_src0_sel_ex),
    .res	(    alu_src0_ex)
);

MUX mux1(
    .src0	(      rf_rd1_ex), 
    .src1	(         imm_ex),
    .sel	(alu_src1_sel_ex),
    .res	(    alu_src1_ex)
);

ALU alu(
    .alu_src0	(    alu_src0_ex), 
    .alu_src1	(    alu_src1_ex),
    .alu_op	(      alu_op_ex),
    .alu_res	(     alu_res_ex)
);

NPC_MUX npc_mux(
    .pc_add4	(      pcadd4_if),
    .pc_offset	(     alu_res_ex),
    .npc_sel	(        npc_sel),
    .npc	(         npc_ex)                
);

Intersegment_REG EX_MEM(
    .clk		(             clk),
    .rst		(             rst),
    .en			(       global_en),
    .stall		(           stall),
    .flush		(            1'b0),
      
    .pcadd4_in		(       pcadd4_ex),
    .pcadd4_out		(      pcadd4_mem),
    .pc_in		(           pc_ex),
    .pc_out		(          pc_mem),
    .inst_in		(         inst_ex),
    .inst_out		(        inst_mem),
    .commit_in		(       commit_ex),
    .commit_out		(      commit_mem),
      
    .imm_in		( 	   imm_ex),
    .imm_out		(         imm_mem),
    .rf_wa_in		(        rf_wa_ex),
    .rf_wa_out		(       rf_wa_mem),
    .rf_rd0_in		(       rf_rd0_ex),
    .rf_rd0_out		(      rf_rd0_mem),
    .rf_rd1_in		(       rf_rd1_ex),
    .rf_rd1_out		(      rf_rd1_mem),
    .rf_we_in		(        rf_we_ex),
    .rf_we_out		(       rf_we_mem),
    .rf_wd_sel_in	(    rf_wd_sel_ex),
    .rf_wd_sel_out	(   rf_wd_sel_mem),
    .alu_op_in		(       alu_op_ex),
    .alu_op_out		(      alu_op_mem),
    .alu_src0_sel_in	( alu_src0_sel_ex),
    .alu_src0_sel_out	(alu_src0_sel_mem),
    .alu_src1_sel_in	( alu_src1_sel_ex),
    .alu_src1_sel_out	(alu_src1_sel_mem),
    .dmem_access_in	(  dmem_access_ex),
    .dmem_access_out	( dmem_access_mem),
    .br_type_in		(      br_type_ex),
    .br_type_out	(     br_type_mem),
    
    .alu_res_in		(      alu_res_ex),
    .alu_res_out	(     alu_res_mem),
            
    .dmem_rd_out_in	(           32'd0),
    .dmem_rd_out_out	(		 ),
    .dmem_wdata_in	(           32'd0),
    .dmem_wdata_out	(	       	 ),
    .dmem_we_in		(      dmem_we_ex),
    .dmem_we_out	(     dmem_we_mem)
);

//for dmem
wire [31 : 0]   dmem_rd_out_mem;
wire [31 : 0]    dmem_rd_out_wb;
wire [31 : 0]    dmem_wdata_mem;
wire [31 : 0]     dmem_wdata_wb;
wire [ 0 : 0]        dmem_we_wb;
assign dmem_addr = alu_res_mem;
assign dmem_wdata = dmem_wdata_mem;
assign dmem_we = dmem_we_mem;

//for MEM/WB
wire [31 : 0]          pcadd4_wb;
wire [31 : 0]              pc_wb;
wire [31 : 0]            inst_wb;
wire [ 0 : 0]          commit_wb;
wire [31 : 0]             imm_wb;
wire [ 4 : 0]           rf_wa_wb;
wire [31 : 0]          rf_rd0_wb;
wire [31 : 0]          rf_rd1_wb;
wire [ 0 : 0]           rf_we_wb;
wire [ 1 : 0]       rf_wd_sel_wb;
wire [ 4 : 0]          alu_op_wb;
wire [ 0 : 0]    alu_src0_sel_wb;
wire [ 0 : 0]    alu_src1_sel_wb;
wire [ 3 : 0]     dmem_access_wb;
wire [ 3 : 0]         br_type_wb;
wire [31 : 0]         alu_res_wb;

SLU slu(
    .addr	(    alu_res_mem),
    .dmem_access(dmem_access_mem),
    .rd_in	(     dmem_rdata),
    .wd_in	(     rf_rd1_mem),
    .rd_out	(dmem_rd_out_mem),
    .wd_out	( dmem_wdata_mem)
);

Intersegment_REG MEM_WB(
    .clk		(             clk),
    .rst		(             rst),
    .en			(       global_en),
    .stall		(           stall),
    .flush		(            1'b0),
      
    .pcadd4_in		(      pcadd4_mem),
    .pcadd4_out		(       pcadd4_wb),
    .pc_in		(          pc_mem),
    .pc_out		(           pc_wb),
    .inst_in		(        inst_mem),
    .inst_out		(         inst_wb),
    .commit_in		(      commit_mem),
    .commit_out		(       commit_wb),
      
    .imm_in		(         imm_mem),
    .imm_out		(          imm_wb),
    .rf_wa_in		(       rf_wa_mem),
    .rf_wa_out		(        rf_wa_wb),
    .rf_rd0_in		(      rf_rd0_mem),
    .rf_rd0_out		(       rf_rd0_wb),
    .rf_rd1_in		(      rf_rd1_mem),
    .rf_rd1_out		(       rf_rd1_wb),
    .rf_we_in		(       rf_we_mem),
    .rf_we_out		(        rf_we_wb),
    .rf_wd_sel_in	(   rf_wd_sel_mem),
    .rf_wd_sel_out	(    rf_wd_sel_wb),
    .alu_op_in		(      alu_op_mem),
    .alu_op_out		(       alu_op_wb),
    .alu_src0_sel_in	(alu_src0_sel_mem),
    .alu_src0_sel_out	( alu_src0_sel_wb),
    .alu_src1_sel_in	(alu_src1_sel_mem),
    .alu_src1_sel_out	( alu_src1_sel_wb),
    .dmem_access_in	( dmem_access_mem),
    .dmem_access_out	(  dmem_access_wb),
    .br_type_in		(     br_type_mem),
    .br_type_out	(      br_type_wb),
    
    .alu_res_in		(     alu_res_mem),
    .alu_res_out	(      alu_res_wb),
            
    .dmem_rd_out_in	( dmem_rd_out_mem),
    .dmem_rd_out_out	(  dmem_rd_out_wb),
    .dmem_wdata_in	(  dmem_wdata_mem),
    .dmem_wdata_out	(   dmem_wdata_wb),
    .dmem_we_in		(     dmem_we_mem),
    .dmem_we_out	(      dmem_we_wb)
);

MUX2 mux2(
    .src0	(     pcadd4_wb), 
    .src1	(    alu_res_wb), 
    .src2	(dmem_rd_out_wb), 
    .src3	(         32'd0),
    .sel	(  rf_wd_sel_wb),
    .res	(      rf_wd_wb)
);

//for commit
reg  [ 0 : 0]   commit_reg          ;
reg  [31 : 0]   commit_pc_reg       ;
reg  [31 : 0]   commit_inst_reg     ;
reg  [ 0 : 0]   commit_halt_reg     ;
reg  [ 0 : 0]   commit_reg_we_reg   ;
reg  [ 4 : 0]   commit_reg_wa_reg   ;
reg  [31 : 0]   commit_reg_wd_reg   ;
reg  [ 0 : 0]   commit_dmem_we_reg  ;
reg  [31 : 0]   commit_dmem_wa_reg  ;
reg  [31 : 0]   commit_dmem_wd_reg  ;

always @(posedge clk) begin
    if (rst) begin
        commit_reg          <= 1'H0;
        commit_pc_reg       <= 32'H0;
        commit_inst_reg     <= 32'H0;
        commit_halt_reg     <= 1'H0;
        commit_reg_we_reg   <= 1'H0;
        commit_reg_wa_reg   <= 5'H0;
        commit_reg_wd_reg   <= 32'H0;
        commit_dmem_we_reg  <= 1'H0;
        commit_dmem_wa_reg  <= 32'H0;
        commit_dmem_wd_reg  <= 32'H0;
    end
    else if (global_en) begin
        commit_reg          <= commit_wb;
        commit_pc_reg       <= pc_wb;
        commit_inst_reg     <= inst_wb;
        commit_halt_reg     <= inst_wb == `HALT_INST;
        commit_reg_we_reg   <= rf_we_wb;
        commit_reg_wa_reg   <= rf_wa_wb;
        commit_reg_wd_reg   <= rf_wd_wb;
        commit_dmem_we_reg  <= dmem_we_wb;                     
        commit_dmem_wa_reg  <= alu_res_wb;                     
        commit_dmem_wd_reg  <= dmem_wdata_wb;                     
    end
end

assign commit               = commit_reg;
assign commit_pc            = commit_pc_reg;
assign commit_inst          = commit_inst_reg;
assign commit_halt          = commit_halt_reg;
assign commit_reg_we        = commit_reg_we_reg;
assign commit_reg_wa        = commit_reg_wa_reg;
assign commit_reg_wd        = commit_reg_wd_reg;
assign commit_dmem_we       = commit_dmem_we_reg;
assign commit_dmem_wa       = commit_dmem_wa_reg;
assign commit_dmem_wd       = commit_dmem_wd_reg;


endmodule


