`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/03/29 18:05:05
// Design Name: 
// Module Name: Adder_LookAhead4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Adder_LookAhead4(
    input [ 3 : 0] a, b,
    input [ 0 : 0] ci, // ���Ե�λ�Ľ�λ
    output [ 3 : 0] s, // ��
    output [ 0 : 0] co // ���λ�Ľ�λ
);

wire [3:0] C;
wire [3:0] G;
wire [3:0] P;
assign G = a & b;
assign P = a ^ b;
assign C[0] = G[0] | ( P[0] & ci );
assign C[1] = G[1] | ( P[1] & G[0] ) | ( P[1] & P[0] & ci );
assign C[2] = G[2] | ( P[2] & G[1] ) | ( P[2] & P[1] & G[0] ) | ( P[2] & P[1] &
P[0] & ci );
assign C[3] = G[3] | ( P[3] & G[2] ) | ( P[3] & P[2] & G[1] ) | ( P[3] & P[2] &
P[1] & G[0] ) | ( P[3] & P[2] & P[1] & P[0] & ci );
assign s[0] = P[0] ^ ci;
assign s[1] = P[1] ^ C[0];
assign s[2] = P[2] ^ C[1];
assign s[3] = P[3] ^ C[2];
assign co = C[3];

endmodule
