
/*
本文件是一个测试文件，用于测试cache模块
工作原理是模仿CPU的读写请求，对cache进行读写操作
将Cache返回的数据与预先数据进行比较，如果一致则测试通过
*/
`timescale 1ns/1ps
module cache_tb();

    //测试参数
    parameter READ_NUM = 2000;  // 测试次数 这里设置为2000次读，1000次写
    parameter WRITE_NUM = 1000;  
    //模块参数
    parameter INDEX_WIDTH       = 3;   // Cache索引位宽 2^3=8行
    parameter LINE_OFFSET_WIDTH = 2;   // 行偏移位宽，决定了一行的宽度 2^2=4字
    parameter SPACE_OFFSET      = 2;   // 一个地址空间占1个字节，因此一个字需要4个地址空间，由于假设为整字读取，处理地址的时候可以默认后两位为0
    parameter MEM_ADDR_WIDTH    = 10;   // 为了简化，这里假设内存地址宽度为10位（CPU请求地址仍然是32位，只不过我们这里简化处理，截断了高位） 
    parameter WAY_NUM           = 1;   // Cache N路组相联(N=1的时候是直接映射)

    // 变化的信号 CPU发出
    reg clk=1;
    reg rstn=1;
    reg stat=0;
    // 等rstn信号稳定后 clk信号才开始翻转
    initial begin
        #1 rstn = 0;
        #1 rstn = 1;
        stat = 1;
    end
    always  #1 clk = ~clk;

    wire [31:0] addr;
    wire r_req;
    wire w_req;
    wire [31:0] w_data;

    // 导线
    wire [31:0] r_data;
    wire miss;
    wire mem_r;
    wire mem_w;
    wire [31:0] mem_addr;
    wire [127:0] mem_w_data;
    wire [127:0] mem_r_data;
    wire mem_ready;

    // 用于测试的信号
    reg [MEM_ADDR_WIDTH-1:0] test_addr[0:READ_NUM+WRITE_NUM-1];  // 用于存储测试地址
    reg [32:0] test_data[0:READ_NUM+WRITE_NUM-1];  // 用于存储测试数据 最高位用于标记是否写入 0：读 1：写
    reg [31:0] test_cnt=0;  // 用于计数，每次读写操作后加1
    reg diff=0;  // 用于标记是否有不一致的数据

    // 用于对比的提交，当前cache应该给出的数据
    wire op;
    wire[31:0] data;
    assign op = test_data[test_cnt-1][32];
    assign data = test_data[test_cnt-1][31:0];
    
    // 状态机
    assign addr = test_addr[test_cnt]<<SPACE_OFFSET;
    assign r_req = test_data[test_cnt][32] == 0 ? 1 : 0;
    assign w_req = test_data[test_cnt][32] == 1 ? 1 : 0;
    assign w_data = test_data[test_cnt][31:0];
    always @(posedge clk) begin
        if (!miss && (test_cnt < READ_NUM+WRITE_NUM) && stat) begin
            if (test_data[test_cnt-1][32] == 0) begin  // 读
                if (r_data != test_data[test_cnt-1][31:0]) begin
                    $display("Read error at %d, expect %h, get %h", test_cnt, test_data[test_cnt-1][31:0], r_data);
                    diff = 1;
                end
            end
            test_cnt <= test_cnt + 1;
        end
    end

    // 例化cache
    cache #(
        .INDEX_WIDTH(INDEX_WIDTH),
        .LINE_OFFSET_WIDTH(LINE_OFFSET_WIDTH),
        .SPACE_OFFSET(SPACE_OFFSET),
        .WAY_NUM(WAY_NUM)
    ) cache_inst(
        .clk(clk),
        .rstn(rstn),
        .addr(addr),
        .r_req(r_req),
        .w_req(w_req),
        .w_data(w_data),
        .r_data(r_data),
        .miss(miss),
        .mem_r(mem_r),
        .mem_w(mem_w),
        .mem_addr(mem_addr),
        .mem_w_data(mem_w_data),
        .mem_r_data(mem_r_data),
        .mem_ready(mem_ready)
    );

    // 内存
    mem #(
        .INDEX_WIDTH(INDEX_WIDTH),
        .LINE_OFFSET_WIDTH(LINE_OFFSET_WIDTH),
        .SPACE_OFFSET(SPACE_OFFSET),
        .MEM_ADDR_WIDTH(MEM_ADDR_WIDTH-LINE_OFFSET_WIDTH),
        .WAY_NUM(WAY_NUM)
    ) mem_inst(
        .clk(clk),
        .rstn(rstn),
        .mem_r(mem_r),
        .mem_w(mem_w),
        .mem_addr(mem_addr),
        .mem_w_data(mem_w_data),
        .mem_r_data(mem_r_data),
        .mem_ready(mem_ready)
    );

    // 初始化测试数据
    initial begin
        test_addr[0] = 0;
        test_data[0] = 33'd2429146761;
        test_addr[1] = 791;
        test_data[1] = 33'd4800218765;
        test_addr[2] = 1;
        test_data[2] = 33'd7700214597;
        test_addr[3] = 2;
        test_data[3] = 33'd244488320;
        test_addr[4] = 337;
        test_data[4] = 33'd2803068549;
        test_addr[5] = 338;
        test_data[5] = 33'd1957293410;
        test_addr[6] = 339;
        test_data[6] = 33'd7213186253;
        test_addr[7] = 340;
        test_data[7] = 33'd3854321255;
        test_addr[8] = 341;
        test_data[8] = 33'd3105826626;
        test_addr[9] = 342;
        test_data[9] = 33'd148146141;
        test_addr[10] = 343;
        test_data[10] = 33'd3938949624;
        test_addr[11] = 344;
        test_data[11] = 33'd477263003;
        test_addr[12] = 345;
        test_data[12] = 33'd7127631255;
        test_addr[13] = 346;
        test_data[13] = 33'd4632375313;
        test_addr[14] = 347;
        test_data[14] = 33'd8330868148;
        test_addr[15] = 348;
        test_data[15] = 33'd3314453200;
        test_addr[16] = 349;
        test_data[16] = 33'd6885446879;
        test_addr[17] = 350;
        test_data[17] = 33'd1842231339;
        test_addr[18] = 351;
        test_data[18] = 33'd8177058853;
        test_addr[19] = 352;
        test_data[19] = 33'd7208142108;
        test_addr[20] = 353;
        test_data[20] = 33'd5225985849;
        test_addr[21] = 354;
        test_data[21] = 33'd369923590;
        test_addr[22] = 355;
        test_data[22] = 33'd2603783369;
        test_addr[23] = 356;
        test_data[23] = 33'd3608961784;
        test_addr[24] = 357;
        test_data[24] = 33'd1704996566;
        test_addr[25] = 358;
        test_data[25] = 33'd3479819972;
        test_addr[26] = 3;
        test_data[26] = 33'd2009627834;
        test_addr[27] = 4;
        test_data[27] = 33'd1187404859;
        test_addr[28] = 5;
        test_data[28] = 33'd7695132375;
        test_addr[29] = 6;
        test_data[29] = 33'd7316665303;
        test_addr[30] = 7;
        test_data[30] = 33'd6930862358;
        test_addr[31] = 8;
        test_data[31] = 33'd4074274575;
        test_addr[32] = 222;
        test_data[32] = 33'd2498690093;
        test_addr[33] = 223;
        test_data[33] = 33'd8269569140;
        test_addr[34] = 224;
        test_data[34] = 33'd4303778506;
        test_addr[35] = 225;
        test_data[35] = 33'd1364845516;
        test_addr[36] = 226;
        test_data[36] = 33'd3088560151;
        test_addr[37] = 227;
        test_data[37] = 33'd4109066461;
        test_addr[38] = 228;
        test_data[38] = 33'd2455014083;
        test_addr[39] = 9;
        test_data[39] = 33'd6453595693;
        test_addr[40] = 10;
        test_data[40] = 33'd2770097472;
        test_addr[41] = 11;
        test_data[41] = 33'd4191856559;
        test_addr[42] = 12;
        test_data[42] = 33'd290304978;
        test_addr[43] = 38;
        test_data[43] = 33'd4009161584;
        test_addr[44] = 39;
        test_data[44] = 33'd2786481955;
        test_addr[45] = 40;
        test_data[45] = 33'd4102836592;
        test_addr[46] = 41;
        test_data[46] = 33'd2145959186;
        test_addr[47] = 42;
        test_data[47] = 33'd527128804;
        test_addr[48] = 43;
        test_data[48] = 33'd3505372607;
        test_addr[49] = 44;
        test_data[49] = 33'd3951540326;
        test_addr[50] = 45;
        test_data[50] = 33'd1124776585;
        test_addr[51] = 46;
        test_data[51] = 33'd1323238552;
        test_addr[52] = 47;
        test_data[52] = 33'd2052202513;
        test_addr[53] = 48;
        test_data[53] = 33'd7512035051;
        test_addr[54] = 49;
        test_data[54] = 33'd8228707208;
        test_addr[55] = 13;
        test_data[55] = 33'd3587268486;
        test_addr[56] = 14;
        test_data[56] = 33'd2853805329;
        test_addr[57] = 15;
        test_data[57] = 33'd7943657238;
        test_addr[58] = 16;
        test_data[58] = 33'd5420650935;
        test_addr[59] = 17;
        test_data[59] = 33'd432400395;
        test_addr[60] = 625;
        test_data[60] = 33'd7533676168;
        test_addr[61] = 626;
        test_data[61] = 33'd4783983235;
        test_addr[62] = 627;
        test_data[62] = 33'd4454129104;
        test_addr[63] = 628;
        test_data[63] = 33'd6593182927;
        test_addr[64] = 629;
        test_data[64] = 33'd1662750713;
        test_addr[65] = 630;
        test_data[65] = 33'd732867767;
        test_addr[66] = 631;
        test_data[66] = 33'd5088069042;
        test_addr[67] = 632;
        test_data[67] = 33'd8427282127;
        test_addr[68] = 633;
        test_data[68] = 33'd3017373220;
        test_addr[69] = 634;
        test_data[69] = 33'd2429702712;
        test_addr[70] = 635;
        test_data[70] = 33'd1607332002;
        test_addr[71] = 636;
        test_data[71] = 33'd6740630795;
        test_addr[72] = 637;
        test_data[72] = 33'd3517993239;
        test_addr[73] = 638;
        test_data[73] = 33'd4136659456;
        test_addr[74] = 639;
        test_data[74] = 33'd86901798;
        test_addr[75] = 640;
        test_data[75] = 33'd3316842311;
        test_addr[76] = 641;
        test_data[76] = 33'd7881353427;
        test_addr[77] = 18;
        test_data[77] = 33'd4089621706;
        test_addr[78] = 19;
        test_data[78] = 33'd2117409300;
        test_addr[79] = 20;
        test_data[79] = 33'd4497406856;
        test_addr[80] = 21;
        test_data[80] = 33'd1866610343;
        test_addr[81] = 22;
        test_data[81] = 33'd5532984872;
        test_addr[82] = 23;
        test_data[82] = 33'd7065585995;
        test_addr[83] = 24;
        test_data[83] = 33'd619906137;
        test_addr[84] = 25;
        test_data[84] = 33'd3881438871;
        test_addr[85] = 26;
        test_data[85] = 33'd1614175349;
        test_addr[86] = 27;
        test_data[86] = 33'd2950000704;
        test_addr[87] = 28;
        test_data[87] = 33'd2040897048;
        test_addr[88] = 29;
        test_data[88] = 33'd580774497;
        test_addr[89] = 30;
        test_data[89] = 33'd7547141517;
        test_addr[90] = 31;
        test_data[90] = 33'd1738403846;
        test_addr[91] = 32;
        test_data[91] = 33'd5133872307;
        test_addr[92] = 33;
        test_data[92] = 33'd5750539502;
        test_addr[93] = 34;
        test_data[93] = 33'd3084178052;
        test_addr[94] = 1011;
        test_data[94] = 33'd4428646174;
        test_addr[95] = 1012;
        test_data[95] = 33'd1486798971;
        test_addr[96] = 1013;
        test_data[96] = 33'd1056707852;
        test_addr[97] = 1014;
        test_data[97] = 33'd414447015;
        test_addr[98] = 1015;
        test_data[98] = 33'd4068782698;
        test_addr[99] = 1016;
        test_data[99] = 33'd379732789;
        test_addr[100] = 1017;
        test_data[100] = 33'd3652225397;
        test_addr[101] = 1018;
        test_data[101] = 33'd2984861369;
        test_addr[102] = 1019;
        test_data[102] = 33'd4093193534;
        test_addr[103] = 1020;
        test_data[103] = 33'd1171431187;
        test_addr[104] = 1021;
        test_data[104] = 33'd4524124189;
        test_addr[105] = 1022;
        test_data[105] = 33'd657762763;
        test_addr[106] = 1023;
        test_data[106] = 33'd2095860060;
        test_addr[107] = 0;
        test_data[107] = 33'd8037811735;
        test_addr[108] = 1;
        test_data[108] = 33'd3405247301;
        test_addr[109] = 2;
        test_data[109] = 33'd244488320;
        test_addr[110] = 3;
        test_data[110] = 33'd2009627834;
        test_addr[111] = 35;
        test_data[111] = 33'd273674846;
        test_addr[112] = 36;
        test_data[112] = 33'd7381012250;
        test_addr[113] = 37;
        test_data[113] = 33'd2005231466;
        test_addr[114] = 38;
        test_data[114] = 33'd4009161584;
        test_addr[115] = 39;
        test_data[115] = 33'd6739391772;
        test_addr[116] = 40;
        test_data[116] = 33'd4962213873;
        test_addr[117] = 41;
        test_data[117] = 33'd5153215001;
        test_addr[118] = 42;
        test_data[118] = 33'd527128804;
        test_addr[119] = 43;
        test_data[119] = 33'd3505372607;
        test_addr[120] = 44;
        test_data[120] = 33'd7703862356;
        test_addr[121] = 45;
        test_data[121] = 33'd1124776585;
        test_addr[122] = 46;
        test_data[122] = 33'd1323238552;
        test_addr[123] = 47;
        test_data[123] = 33'd4462151347;
        test_addr[124] = 48;
        test_data[124] = 33'd3217067755;
        test_addr[125] = 49;
        test_data[125] = 33'd3933739912;
        test_addr[126] = 50;
        test_data[126] = 33'd7124950387;
        test_addr[127] = 1008;
        test_data[127] = 33'd4215858546;
        test_addr[128] = 1009;
        test_data[128] = 33'd1316389492;
        test_addr[129] = 1010;
        test_data[129] = 33'd3511528593;
        test_addr[130] = 1011;
        test_data[130] = 33'd133678878;
        test_addr[131] = 1012;
        test_data[131] = 33'd1486798971;
        test_addr[132] = 1013;
        test_data[132] = 33'd1056707852;
        test_addr[133] = 51;
        test_data[133] = 33'd2194417863;
        test_addr[134] = 52;
        test_data[134] = 33'd4539344385;
        test_addr[135] = 53;
        test_data[135] = 33'd1748677916;
        test_addr[136] = 989;
        test_data[136] = 33'd3635546882;
        test_addr[137] = 990;
        test_data[137] = 33'd7674610783;
        test_addr[138] = 991;
        test_data[138] = 33'd5407353489;
        test_addr[139] = 992;
        test_data[139] = 33'd5259146489;
        test_addr[140] = 993;
        test_data[140] = 33'd1857244546;
        test_addr[141] = 54;
        test_data[141] = 33'd2532063245;
        test_addr[142] = 55;
        test_data[142] = 33'd2155416609;
        test_addr[143] = 56;
        test_data[143] = 33'd2965160517;
        test_addr[144] = 57;
        test_data[144] = 33'd4360448829;
        test_addr[145] = 58;
        test_data[145] = 33'd3980185017;
        test_addr[146] = 13;
        test_data[146] = 33'd3587268486;
        test_addr[147] = 14;
        test_data[147] = 33'd5473352741;
        test_addr[148] = 15;
        test_data[148] = 33'd3648689942;
        test_addr[149] = 16;
        test_data[149] = 33'd1125683639;
        test_addr[150] = 17;
        test_data[150] = 33'd4435668262;
        test_addr[151] = 18;
        test_data[151] = 33'd4089621706;
        test_addr[152] = 19;
        test_data[152] = 33'd6905529021;
        test_addr[153] = 20;
        test_data[153] = 33'd6214605454;
        test_addr[154] = 21;
        test_data[154] = 33'd1866610343;
        test_addr[155] = 22;
        test_data[155] = 33'd1238017576;
        test_addr[156] = 23;
        test_data[156] = 33'd2770618699;
        test_addr[157] = 59;
        test_data[157] = 33'd587109440;
        test_addr[158] = 60;
        test_data[158] = 33'd2464752507;
        test_addr[159] = 61;
        test_data[159] = 33'd3065752321;
        test_addr[160] = 62;
        test_data[160] = 33'd3712003529;
        test_addr[161] = 63;
        test_data[161] = 33'd807961889;
        test_addr[162] = 54;
        test_data[162] = 33'd2532063245;
        test_addr[163] = 55;
        test_data[163] = 33'd2155416609;
        test_addr[164] = 56;
        test_data[164] = 33'd2965160517;
        test_addr[165] = 57;
        test_data[165] = 33'd65481533;
        test_addr[166] = 58;
        test_data[166] = 33'd3980185017;
        test_addr[167] = 59;
        test_data[167] = 33'd587109440;
        test_addr[168] = 60;
        test_data[168] = 33'd2464752507;
        test_addr[169] = 61;
        test_data[169] = 33'd3065752321;
        test_addr[170] = 62;
        test_data[170] = 33'd3712003529;
        test_addr[171] = 64;
        test_data[171] = 33'd7302595289;
        test_addr[172] = 65;
        test_data[172] = 33'd1673314307;
        test_addr[173] = 66;
        test_data[173] = 33'd5228628;
        test_addr[174] = 67;
        test_data[174] = 33'd283800910;
        test_addr[175] = 68;
        test_data[175] = 33'd3879425881;
        test_addr[176] = 69;
        test_data[176] = 33'd2408633668;
        test_addr[177] = 70;
        test_data[177] = 33'd6358267530;
        test_addr[178] = 71;
        test_data[178] = 33'd3398690954;
        test_addr[179] = 72;
        test_data[179] = 33'd583387573;
        test_addr[180] = 73;
        test_data[180] = 33'd1855683855;
        test_addr[181] = 74;
        test_data[181] = 33'd1226571034;
        test_addr[182] = 75;
        test_data[182] = 33'd1317445743;
        test_addr[183] = 76;
        test_data[183] = 33'd2183571412;
        test_addr[184] = 291;
        test_data[184] = 33'd7426318834;
        test_addr[185] = 292;
        test_data[185] = 33'd149615558;
        test_addr[186] = 293;
        test_data[186] = 33'd880389596;
        test_addr[187] = 294;
        test_data[187] = 33'd6791871258;
        test_addr[188] = 295;
        test_data[188] = 33'd1453477040;
        test_addr[189] = 296;
        test_data[189] = 33'd72603561;
        test_addr[190] = 297;
        test_data[190] = 33'd6067958687;
        test_addr[191] = 77;
        test_data[191] = 33'd1951277074;
        test_addr[192] = 827;
        test_data[192] = 33'd4087048189;
        test_addr[193] = 828;
        test_data[193] = 33'd3346872234;
        test_addr[194] = 829;
        test_data[194] = 33'd275433189;
        test_addr[195] = 830;
        test_data[195] = 33'd3958563769;
        test_addr[196] = 831;
        test_data[196] = 33'd6074066124;
        test_addr[197] = 832;
        test_data[197] = 33'd2891161115;
        test_addr[198] = 833;
        test_data[198] = 33'd1793456890;
        test_addr[199] = 834;
        test_data[199] = 33'd3031697508;
        test_addr[200] = 835;
        test_data[200] = 33'd6861685134;
        test_addr[201] = 836;
        test_data[201] = 33'd319479514;
        test_addr[202] = 837;
        test_data[202] = 33'd6856140373;
        test_addr[203] = 838;
        test_data[203] = 33'd2155428742;
        test_addr[204] = 839;
        test_data[204] = 33'd2174987116;
        test_addr[205] = 840;
        test_data[205] = 33'd403783328;
        test_addr[206] = 841;
        test_data[206] = 33'd846659615;
        test_addr[207] = 78;
        test_data[207] = 33'd3938077862;
        test_addr[208] = 79;
        test_data[208] = 33'd3352086201;
        test_addr[209] = 80;
        test_data[209] = 33'd5635362666;
        test_addr[210] = 81;
        test_data[210] = 33'd7615811479;
        test_addr[211] = 82;
        test_data[211] = 33'd2763428529;
        test_addr[212] = 963;
        test_data[212] = 33'd3778906056;
        test_addr[213] = 964;
        test_data[213] = 33'd1676243570;
        test_addr[214] = 965;
        test_data[214] = 33'd533232901;
        test_addr[215] = 966;
        test_data[215] = 33'd168242151;
        test_addr[216] = 967;
        test_data[216] = 33'd2540554632;
        test_addr[217] = 968;
        test_data[217] = 33'd759450314;
        test_addr[218] = 969;
        test_data[218] = 33'd4246657183;
        test_addr[219] = 970;
        test_data[219] = 33'd1523162636;
        test_addr[220] = 971;
        test_data[220] = 33'd1160760996;
        test_addr[221] = 972;
        test_data[221] = 33'd764522856;
        test_addr[222] = 973;
        test_data[222] = 33'd1572552106;
        test_addr[223] = 974;
        test_data[223] = 33'd3026688618;
        test_addr[224] = 975;
        test_data[224] = 33'd902628290;
        test_addr[225] = 976;
        test_data[225] = 33'd7246384212;
        test_addr[226] = 977;
        test_data[226] = 33'd275231142;
        test_addr[227] = 978;
        test_data[227] = 33'd6633914448;
        test_addr[228] = 979;
        test_data[228] = 33'd2852800281;
        test_addr[229] = 980;
        test_data[229] = 33'd2034359482;
        test_addr[230] = 981;
        test_data[230] = 33'd4613200403;
        test_addr[231] = 83;
        test_data[231] = 33'd1828590022;
        test_addr[232] = 84;
        test_data[232] = 33'd1081301073;
        test_addr[233] = 655;
        test_data[233] = 33'd4383732844;
        test_addr[234] = 656;
        test_data[234] = 33'd2492457321;
        test_addr[235] = 657;
        test_data[235] = 33'd576451002;
        test_addr[236] = 658;
        test_data[236] = 33'd4466531428;
        test_addr[237] = 659;
        test_data[237] = 33'd4136402978;
        test_addr[238] = 660;
        test_data[238] = 33'd6452148123;
        test_addr[239] = 661;
        test_data[239] = 33'd1404351648;
        test_addr[240] = 662;
        test_data[240] = 33'd4126887004;
        test_addr[241] = 663;
        test_data[241] = 33'd3355262986;
        test_addr[242] = 664;
        test_data[242] = 33'd1318050398;
        test_addr[243] = 665;
        test_data[243] = 33'd5293634356;
        test_addr[244] = 666;
        test_data[244] = 33'd8340347185;
        test_addr[245] = 667;
        test_data[245] = 33'd1268036190;
        test_addr[246] = 668;
        test_data[246] = 33'd5869128725;
        test_addr[247] = 669;
        test_data[247] = 33'd7667091059;
        test_addr[248] = 670;
        test_data[248] = 33'd2901628700;
        test_addr[249] = 671;
        test_data[249] = 33'd3009182528;
        test_addr[250] = 672;
        test_data[250] = 33'd7649982545;
        test_addr[251] = 673;
        test_data[251] = 33'd3204904385;
        test_addr[252] = 674;
        test_data[252] = 33'd6685950640;
        test_addr[253] = 675;
        test_data[253] = 33'd2709261325;
        test_addr[254] = 676;
        test_data[254] = 33'd1104785019;
        test_addr[255] = 677;
        test_data[255] = 33'd1594126675;
        test_addr[256] = 678;
        test_data[256] = 33'd4257693411;
        test_addr[257] = 679;
        test_data[257] = 33'd4395771824;
        test_addr[258] = 680;
        test_data[258] = 33'd7414008368;
        test_addr[259] = 681;
        test_data[259] = 33'd1236016341;
        test_addr[260] = 682;
        test_data[260] = 33'd6984815728;
        test_addr[261] = 683;
        test_data[261] = 33'd3097106317;
        test_addr[262] = 85;
        test_data[262] = 33'd725363894;
        test_addr[263] = 86;
        test_data[263] = 33'd1595499640;
        test_addr[264] = 87;
        test_data[264] = 33'd597900638;
        test_addr[265] = 88;
        test_data[265] = 33'd1179514588;
        test_addr[266] = 89;
        test_data[266] = 33'd4756071467;
        test_addr[267] = 90;
        test_data[267] = 33'd43380869;
        test_addr[268] = 91;
        test_data[268] = 33'd138001890;
        test_addr[269] = 92;
        test_data[269] = 33'd403469968;
        test_addr[270] = 93;
        test_data[270] = 33'd563973034;
        test_addr[271] = 94;
        test_data[271] = 33'd8508161183;
        test_addr[272] = 95;
        test_data[272] = 33'd610452162;
        test_addr[273] = 96;
        test_data[273] = 33'd2080744587;
        test_addr[274] = 97;
        test_data[274] = 33'd654962339;
        test_addr[275] = 98;
        test_data[275] = 33'd3684430035;
        test_addr[276] = 99;
        test_data[276] = 33'd1718939551;
        test_addr[277] = 100;
        test_data[277] = 33'd3845605637;
        test_addr[278] = 101;
        test_data[278] = 33'd669798772;
        test_addr[279] = 102;
        test_data[279] = 33'd746597445;
        test_addr[280] = 103;
        test_data[280] = 33'd5454673078;
        test_addr[281] = 104;
        test_data[281] = 33'd7617652761;
        test_addr[282] = 105;
        test_data[282] = 33'd1511183284;
        test_addr[283] = 106;
        test_data[283] = 33'd1630641212;
        test_addr[284] = 107;
        test_data[284] = 33'd4002934247;
        test_addr[285] = 108;
        test_data[285] = 33'd5424746931;
        test_addr[286] = 109;
        test_data[286] = 33'd1300879613;
        test_addr[287] = 110;
        test_data[287] = 33'd1563193765;
        test_addr[288] = 111;
        test_data[288] = 33'd59269632;
        test_addr[289] = 112;
        test_data[289] = 33'd26118987;
        test_addr[290] = 113;
        test_data[290] = 33'd124869335;
        test_addr[291] = 114;
        test_data[291] = 33'd4558599183;
        test_addr[292] = 710;
        test_data[292] = 33'd3654683160;
        test_addr[293] = 711;
        test_data[293] = 33'd1104666845;
        test_addr[294] = 712;
        test_data[294] = 33'd3993640537;
        test_addr[295] = 713;
        test_data[295] = 33'd3877347980;
        test_addr[296] = 714;
        test_data[296] = 33'd1793666688;
        test_addr[297] = 115;
        test_data[297] = 33'd2227853741;
        test_addr[298] = 116;
        test_data[298] = 33'd6428178809;
        test_addr[299] = 117;
        test_data[299] = 33'd5778825445;
        test_addr[300] = 118;
        test_data[300] = 33'd2838500611;
        test_addr[301] = 119;
        test_data[301] = 33'd8190291852;
        test_addr[302] = 120;
        test_data[302] = 33'd5300811407;
        test_addr[303] = 121;
        test_data[303] = 33'd539709361;
        test_addr[304] = 51;
        test_data[304] = 33'd2194417863;
        test_addr[305] = 52;
        test_data[305] = 33'd244377089;
        test_addr[306] = 53;
        test_data[306] = 33'd1748677916;
        test_addr[307] = 54;
        test_data[307] = 33'd8327263198;
        test_addr[308] = 122;
        test_data[308] = 33'd3741684855;
        test_addr[309] = 123;
        test_data[309] = 33'd2458661410;
        test_addr[310] = 124;
        test_data[310] = 33'd7156413009;
        test_addr[311] = 125;
        test_data[311] = 33'd5171785345;
        test_addr[312] = 126;
        test_data[312] = 33'd4195730453;
        test_addr[313] = 592;
        test_data[313] = 33'd3656952568;
        test_addr[314] = 593;
        test_data[314] = 33'd767211102;
        test_addr[315] = 127;
        test_data[315] = 33'd4971126949;
        test_addr[316] = 128;
        test_data[316] = 33'd6055166934;
        test_addr[317] = 129;
        test_data[317] = 33'd652071928;
        test_addr[318] = 130;
        test_data[318] = 33'd4776256812;
        test_addr[319] = 131;
        test_data[319] = 33'd6515894620;
        test_addr[320] = 132;
        test_data[320] = 33'd3352808087;
        test_addr[321] = 133;
        test_data[321] = 33'd2182795532;
        test_addr[322] = 134;
        test_data[322] = 33'd7198008121;
        test_addr[323] = 135;
        test_data[323] = 33'd2176215843;
        test_addr[324] = 136;
        test_data[324] = 33'd3446836288;
        test_addr[325] = 137;
        test_data[325] = 33'd2464351703;
        test_addr[326] = 138;
        test_data[326] = 33'd8552288077;
        test_addr[327] = 139;
        test_data[327] = 33'd7895743433;
        test_addr[328] = 140;
        test_data[328] = 33'd3314446855;
        test_addr[329] = 141;
        test_data[329] = 33'd1108123326;
        test_addr[330] = 142;
        test_data[330] = 33'd6820992057;
        test_addr[331] = 986;
        test_data[331] = 33'd1388652941;
        test_addr[332] = 987;
        test_data[332] = 33'd7332995067;
        test_addr[333] = 988;
        test_data[333] = 33'd2478676154;
        test_addr[334] = 989;
        test_data[334] = 33'd3635546882;
        test_addr[335] = 990;
        test_data[335] = 33'd3379643487;
        test_addr[336] = 991;
        test_data[336] = 33'd1112386193;
        test_addr[337] = 992;
        test_data[337] = 33'd964179193;
        test_addr[338] = 993;
        test_data[338] = 33'd1857244546;
        test_addr[339] = 994;
        test_data[339] = 33'd2089204886;
        test_addr[340] = 995;
        test_data[340] = 33'd3226654615;
        test_addr[341] = 996;
        test_data[341] = 33'd3922015050;
        test_addr[342] = 997;
        test_data[342] = 33'd1759334156;
        test_addr[343] = 998;
        test_data[343] = 33'd6923401218;
        test_addr[344] = 999;
        test_data[344] = 33'd3093736890;
        test_addr[345] = 1000;
        test_data[345] = 33'd4411027836;
        test_addr[346] = 143;
        test_data[346] = 33'd1862437858;
        test_addr[347] = 144;
        test_data[347] = 33'd8371171917;
        test_addr[348] = 145;
        test_data[348] = 33'd5906598566;
        test_addr[349] = 540;
        test_data[349] = 33'd4853221104;
        test_addr[350] = 541;
        test_data[350] = 33'd1920105602;
        test_addr[351] = 542;
        test_data[351] = 33'd3693452330;
        test_addr[352] = 543;
        test_data[352] = 33'd6226430920;
        test_addr[353] = 544;
        test_data[353] = 33'd118999468;
        test_addr[354] = 545;
        test_data[354] = 33'd1749290836;
        test_addr[355] = 546;
        test_data[355] = 33'd717909476;
        test_addr[356] = 547;
        test_data[356] = 33'd1656097789;
        test_addr[357] = 548;
        test_data[357] = 33'd3975122350;
        test_addr[358] = 549;
        test_data[358] = 33'd2127589844;
        test_addr[359] = 550;
        test_data[359] = 33'd7673183117;
        test_addr[360] = 551;
        test_data[360] = 33'd7845091920;
        test_addr[361] = 552;
        test_data[361] = 33'd1286678884;
        test_addr[362] = 553;
        test_data[362] = 33'd1687299562;
        test_addr[363] = 554;
        test_data[363] = 33'd3923557028;
        test_addr[364] = 555;
        test_data[364] = 33'd2248499919;
        test_addr[365] = 556;
        test_data[365] = 33'd2939472687;
        test_addr[366] = 557;
        test_data[366] = 33'd985122537;
        test_addr[367] = 558;
        test_data[367] = 33'd3808977718;
        test_addr[368] = 559;
        test_data[368] = 33'd839457297;
        test_addr[369] = 560;
        test_data[369] = 33'd7254175320;
        test_addr[370] = 561;
        test_data[370] = 33'd5112667199;
        test_addr[371] = 146;
        test_data[371] = 33'd3958907471;
        test_addr[372] = 147;
        test_data[372] = 33'd3396137010;
        test_addr[373] = 148;
        test_data[373] = 33'd5621973513;
        test_addr[374] = 149;
        test_data[374] = 33'd5771382092;
        test_addr[375] = 150;
        test_data[375] = 33'd2726814038;
        test_addr[376] = 151;
        test_data[376] = 33'd4527197915;
        test_addr[377] = 152;
        test_data[377] = 33'd800774714;
        test_addr[378] = 153;
        test_data[378] = 33'd7642976212;
        test_addr[379] = 154;
        test_data[379] = 33'd3022540257;
        test_addr[380] = 155;
        test_data[380] = 33'd5928842315;
        test_addr[381] = 156;
        test_data[381] = 33'd5292043467;
        test_addr[382] = 157;
        test_data[382] = 33'd98365346;
        test_addr[383] = 158;
        test_data[383] = 33'd2430407245;
        test_addr[384] = 159;
        test_data[384] = 33'd5170958586;
        test_addr[385] = 160;
        test_data[385] = 33'd2802001540;
        test_addr[386] = 161;
        test_data[386] = 33'd260760954;
        test_addr[387] = 162;
        test_data[387] = 33'd760186910;
        test_addr[388] = 291;
        test_data[388] = 33'd3131351538;
        test_addr[389] = 292;
        test_data[389] = 33'd149615558;
        test_addr[390] = 293;
        test_data[390] = 33'd880389596;
        test_addr[391] = 294;
        test_data[391] = 33'd8360622715;
        test_addr[392] = 295;
        test_data[392] = 33'd1453477040;
        test_addr[393] = 163;
        test_data[393] = 33'd2417096706;
        test_addr[394] = 164;
        test_data[394] = 33'd3847429411;
        test_addr[395] = 165;
        test_data[395] = 33'd7228023884;
        test_addr[396] = 166;
        test_data[396] = 33'd1567391663;
        test_addr[397] = 326;
        test_data[397] = 33'd7506007486;
        test_addr[398] = 327;
        test_data[398] = 33'd4021375997;
        test_addr[399] = 328;
        test_data[399] = 33'd4211559137;
        test_addr[400] = 329;
        test_data[400] = 33'd508970632;
        test_addr[401] = 330;
        test_data[401] = 33'd2871069657;
        test_addr[402] = 331;
        test_data[402] = 33'd7316552142;
        test_addr[403] = 332;
        test_data[403] = 33'd8097508361;
        test_addr[404] = 333;
        test_data[404] = 33'd3777587601;
        test_addr[405] = 334;
        test_data[405] = 33'd2560750633;
        test_addr[406] = 167;
        test_data[406] = 33'd4201079425;
        test_addr[407] = 821;
        test_data[407] = 33'd3918583867;
        test_addr[408] = 822;
        test_data[408] = 33'd3241601505;
        test_addr[409] = 823;
        test_data[409] = 33'd3228310104;
        test_addr[410] = 824;
        test_data[410] = 33'd1705558585;
        test_addr[411] = 825;
        test_data[411] = 33'd3901277367;
        test_addr[412] = 826;
        test_data[412] = 33'd4536649406;
        test_addr[413] = 827;
        test_data[413] = 33'd6028813588;
        test_addr[414] = 828;
        test_data[414] = 33'd3346872234;
        test_addr[415] = 829;
        test_data[415] = 33'd5963846806;
        test_addr[416] = 830;
        test_data[416] = 33'd3958563769;
        test_addr[417] = 831;
        test_data[417] = 33'd5911680679;
        test_addr[418] = 832;
        test_data[418] = 33'd2891161115;
        test_addr[419] = 833;
        test_data[419] = 33'd5517701565;
        test_addr[420] = 834;
        test_data[420] = 33'd3031697508;
        test_addr[421] = 835;
        test_data[421] = 33'd2566717838;
        test_addr[422] = 836;
        test_data[422] = 33'd4874452461;
        test_addr[423] = 837;
        test_data[423] = 33'd2561173077;
        test_addr[424] = 838;
        test_data[424] = 33'd6744048819;
        test_addr[425] = 168;
        test_data[425] = 33'd244697080;
        test_addr[426] = 169;
        test_data[426] = 33'd5768117693;
        test_addr[427] = 170;
        test_data[427] = 33'd6007450025;
        test_addr[428] = 171;
        test_data[428] = 33'd4446887705;
        test_addr[429] = 172;
        test_data[429] = 33'd2706684257;
        test_addr[430] = 173;
        test_data[430] = 33'd1739717906;
        test_addr[431] = 174;
        test_data[431] = 33'd8319474124;
        test_addr[432] = 175;
        test_data[432] = 33'd1951074742;
        test_addr[433] = 176;
        test_data[433] = 33'd3605693122;
        test_addr[434] = 177;
        test_data[434] = 33'd6842266167;
        test_addr[435] = 178;
        test_data[435] = 33'd1390194371;
        test_addr[436] = 179;
        test_data[436] = 33'd4169806564;
        test_addr[437] = 180;
        test_data[437] = 33'd2888358889;
        test_addr[438] = 181;
        test_data[438] = 33'd485480945;
        test_addr[439] = 182;
        test_data[439] = 33'd407882722;
        test_addr[440] = 183;
        test_data[440] = 33'd1700753432;
        test_addr[441] = 184;
        test_data[441] = 33'd4125218622;
        test_addr[442] = 185;
        test_data[442] = 33'd5140063103;
        test_addr[443] = 186;
        test_data[443] = 33'd621023615;
        test_addr[444] = 187;
        test_data[444] = 33'd4624618666;
        test_addr[445] = 188;
        test_data[445] = 33'd3828919794;
        test_addr[446] = 189;
        test_data[446] = 33'd2152553771;
        test_addr[447] = 190;
        test_data[447] = 33'd2871768144;
        test_addr[448] = 456;
        test_data[448] = 33'd2655493248;
        test_addr[449] = 457;
        test_data[449] = 33'd2493953492;
        test_addr[450] = 458;
        test_data[450] = 33'd2786993620;
        test_addr[451] = 459;
        test_data[451] = 33'd5121202977;
        test_addr[452] = 460;
        test_data[452] = 33'd7685281244;
        test_addr[453] = 461;
        test_data[453] = 33'd5915799328;
        test_addr[454] = 462;
        test_data[454] = 33'd8065079457;
        test_addr[455] = 463;
        test_data[455] = 33'd2623477901;
        test_addr[456] = 464;
        test_data[456] = 33'd7442112983;
        test_addr[457] = 465;
        test_data[457] = 33'd6345593786;
        test_addr[458] = 466;
        test_data[458] = 33'd3459645207;
        test_addr[459] = 467;
        test_data[459] = 33'd6832024842;
        test_addr[460] = 468;
        test_data[460] = 33'd3992930714;
        test_addr[461] = 469;
        test_data[461] = 33'd1664670904;
        test_addr[462] = 470;
        test_data[462] = 33'd7559203245;
        test_addr[463] = 471;
        test_data[463] = 33'd4727862512;
        test_addr[464] = 472;
        test_data[464] = 33'd8487967563;
        test_addr[465] = 473;
        test_data[465] = 33'd1293966191;
        test_addr[466] = 474;
        test_data[466] = 33'd8003696540;
        test_addr[467] = 475;
        test_data[467] = 33'd2268014519;
        test_addr[468] = 476;
        test_data[468] = 33'd3560019982;
        test_addr[469] = 477;
        test_data[469] = 33'd3221152013;
        test_addr[470] = 478;
        test_data[470] = 33'd5522729664;
        test_addr[471] = 479;
        test_data[471] = 33'd2603322669;
        test_addr[472] = 191;
        test_data[472] = 33'd5954101850;
        test_addr[473] = 192;
        test_data[473] = 33'd4618404879;
        test_addr[474] = 193;
        test_data[474] = 33'd1908158991;
        test_addr[475] = 194;
        test_data[475] = 33'd3455513250;
        test_addr[476] = 195;
        test_data[476] = 33'd7314517096;
        test_addr[477] = 196;
        test_data[477] = 33'd3889204301;
        test_addr[478] = 197;
        test_data[478] = 33'd3675913621;
        test_addr[479] = 198;
        test_data[479] = 33'd400801465;
        test_addr[480] = 199;
        test_data[480] = 33'd8286985878;
        test_addr[481] = 200;
        test_data[481] = 33'd3223549335;
        test_addr[482] = 201;
        test_data[482] = 33'd2012336102;
        test_addr[483] = 491;
        test_data[483] = 33'd6404490069;
        test_addr[484] = 492;
        test_data[484] = 33'd712901222;
        test_addr[485] = 493;
        test_data[485] = 33'd712725379;
        test_addr[486] = 494;
        test_data[486] = 33'd4592674516;
        test_addr[487] = 202;
        test_data[487] = 33'd631181234;
        test_addr[488] = 203;
        test_data[488] = 33'd6980300848;
        test_addr[489] = 204;
        test_data[489] = 33'd7522611158;
        test_addr[490] = 205;
        test_data[490] = 33'd540360476;
        test_addr[491] = 43;
        test_data[491] = 33'd6061199720;
        test_addr[492] = 44;
        test_data[492] = 33'd7824797516;
        test_addr[493] = 45;
        test_data[493] = 33'd1124776585;
        test_addr[494] = 206;
        test_data[494] = 33'd2946247101;
        test_addr[495] = 207;
        test_data[495] = 33'd689273551;
        test_addr[496] = 208;
        test_data[496] = 33'd1843892378;
        test_addr[497] = 209;
        test_data[497] = 33'd6979028179;
        test_addr[498] = 210;
        test_data[498] = 33'd4727038944;
        test_addr[499] = 211;
        test_data[499] = 33'd3948687695;
        test_addr[500] = 695;
        test_data[500] = 33'd4120276502;
        test_addr[501] = 696;
        test_data[501] = 33'd1053390424;
        test_addr[502] = 697;
        test_data[502] = 33'd6590853502;
        test_addr[503] = 698;
        test_data[503] = 33'd5270229509;
        test_addr[504] = 699;
        test_data[504] = 33'd7268085778;
        test_addr[505] = 700;
        test_data[505] = 33'd5263355905;
        test_addr[506] = 701;
        test_data[506] = 33'd835744670;
        test_addr[507] = 702;
        test_data[507] = 33'd3588029089;
        test_addr[508] = 703;
        test_data[508] = 33'd1255659046;
        test_addr[509] = 704;
        test_data[509] = 33'd998116682;
        test_addr[510] = 705;
        test_data[510] = 33'd6206225240;
        test_addr[511] = 706;
        test_data[511] = 33'd7816345375;
        test_addr[512] = 212;
        test_data[512] = 33'd8192542853;
        test_addr[513] = 213;
        test_data[513] = 33'd6157732905;
        test_addr[514] = 214;
        test_data[514] = 33'd3563881117;
        test_addr[515] = 215;
        test_data[515] = 33'd4879403786;
        test_addr[516] = 242;
        test_data[516] = 33'd8114562116;
        test_addr[517] = 243;
        test_data[517] = 33'd309132402;
        test_addr[518] = 244;
        test_data[518] = 33'd3986444448;
        test_addr[519] = 245;
        test_data[519] = 33'd7804312792;
        test_addr[520] = 246;
        test_data[520] = 33'd2440705799;
        test_addr[521] = 247;
        test_data[521] = 33'd7052191550;
        test_addr[522] = 248;
        test_data[522] = 33'd1851737756;
        test_addr[523] = 249;
        test_data[523] = 33'd4121500431;
        test_addr[524] = 250;
        test_data[524] = 33'd1892908102;
        test_addr[525] = 251;
        test_data[525] = 33'd4348416482;
        test_addr[526] = 252;
        test_data[526] = 33'd4633393528;
        test_addr[527] = 253;
        test_data[527] = 33'd1046892784;
        test_addr[528] = 254;
        test_data[528] = 33'd893686890;
        test_addr[529] = 255;
        test_data[529] = 33'd738701221;
        test_addr[530] = 256;
        test_data[530] = 33'd104124540;
        test_addr[531] = 257;
        test_data[531] = 33'd2272834637;
        test_addr[532] = 258;
        test_data[532] = 33'd7413699645;
        test_addr[533] = 259;
        test_data[533] = 33'd3199409289;
        test_addr[534] = 260;
        test_data[534] = 33'd3784376997;
        test_addr[535] = 261;
        test_data[535] = 33'd3435254937;
        test_addr[536] = 262;
        test_data[536] = 33'd7488855415;
        test_addr[537] = 263;
        test_data[537] = 33'd1168259603;
        test_addr[538] = 264;
        test_data[538] = 33'd3017312274;
        test_addr[539] = 265;
        test_data[539] = 33'd4232753553;
        test_addr[540] = 266;
        test_data[540] = 33'd4193755358;
        test_addr[541] = 267;
        test_data[541] = 33'd2420869187;
        test_addr[542] = 268;
        test_data[542] = 33'd2644833872;
        test_addr[543] = 269;
        test_data[543] = 33'd2018394395;
        test_addr[544] = 270;
        test_data[544] = 33'd6329395444;
        test_addr[545] = 271;
        test_data[545] = 33'd4226387963;
        test_addr[546] = 272;
        test_data[546] = 33'd1785668236;
        test_addr[547] = 273;
        test_data[547] = 33'd7147254911;
        test_addr[548] = 274;
        test_data[548] = 33'd3297475855;
        test_addr[549] = 275;
        test_data[549] = 33'd4315669401;
        test_addr[550] = 276;
        test_data[550] = 33'd151084863;
        test_addr[551] = 277;
        test_data[551] = 33'd1313409944;
        test_addr[552] = 278;
        test_data[552] = 33'd3951155712;
        test_addr[553] = 279;
        test_data[553] = 33'd2152272633;
        test_addr[554] = 280;
        test_data[554] = 33'd1318904363;
        test_addr[555] = 281;
        test_data[555] = 33'd5814186882;
        test_addr[556] = 282;
        test_data[556] = 33'd4737997644;
        test_addr[557] = 283;
        test_data[557] = 33'd1573656911;
        test_addr[558] = 284;
        test_data[558] = 33'd8111976187;
        test_addr[559] = 285;
        test_data[559] = 33'd8373853213;
        test_addr[560] = 216;
        test_data[560] = 33'd313568208;
        test_addr[561] = 389;
        test_data[561] = 33'd6538596791;
        test_addr[562] = 217;
        test_data[562] = 33'd6468322402;
        test_addr[563] = 488;
        test_data[563] = 33'd3725295247;
        test_addr[564] = 489;
        test_data[564] = 33'd2421545610;
        test_addr[565] = 490;
        test_data[565] = 33'd3475954419;
        test_addr[566] = 491;
        test_data[566] = 33'd2109522773;
        test_addr[567] = 492;
        test_data[567] = 33'd712901222;
        test_addr[568] = 493;
        test_data[568] = 33'd712725379;
        test_addr[569] = 494;
        test_data[569] = 33'd297707220;
        test_addr[570] = 495;
        test_data[570] = 33'd5054457440;
        test_addr[571] = 496;
        test_data[571] = 33'd822810503;
        test_addr[572] = 497;
        test_data[572] = 33'd1711199328;
        test_addr[573] = 498;
        test_data[573] = 33'd3738045385;
        test_addr[574] = 499;
        test_data[574] = 33'd3460457963;
        test_addr[575] = 500;
        test_data[575] = 33'd4507997725;
        test_addr[576] = 501;
        test_data[576] = 33'd6104803262;
        test_addr[577] = 502;
        test_data[577] = 33'd2391045745;
        test_addr[578] = 218;
        test_data[578] = 33'd3295815568;
        test_addr[579] = 219;
        test_data[579] = 33'd1970268263;
        test_addr[580] = 220;
        test_data[580] = 33'd3319839920;
        test_addr[581] = 221;
        test_data[581] = 33'd2679756236;
        test_addr[582] = 222;
        test_data[582] = 33'd2498690093;
        test_addr[583] = 223;
        test_data[583] = 33'd3974601844;
        test_addr[584] = 224;
        test_data[584] = 33'd8811210;
        test_addr[585] = 225;
        test_data[585] = 33'd7519316143;
        test_addr[586] = 226;
        test_data[586] = 33'd6726459389;
        test_addr[587] = 227;
        test_data[587] = 33'd4109066461;
        test_addr[588] = 228;
        test_data[588] = 33'd7322327114;
        test_addr[589] = 646;
        test_data[589] = 33'd1560612810;
        test_addr[590] = 647;
        test_data[590] = 33'd360683726;
        test_addr[591] = 648;
        test_data[591] = 33'd2360713956;
        test_addr[592] = 649;
        test_data[592] = 33'd7644754019;
        test_addr[593] = 650;
        test_data[593] = 33'd4203221935;
        test_addr[594] = 229;
        test_data[594] = 33'd2383148880;
        test_addr[595] = 984;
        test_data[595] = 33'd7137525381;
        test_addr[596] = 985;
        test_data[596] = 33'd1224700992;
        test_addr[597] = 986;
        test_data[597] = 33'd5821328108;
        test_addr[598] = 987;
        test_data[598] = 33'd3038027771;
        test_addr[599] = 988;
        test_data[599] = 33'd4566854779;
        test_addr[600] = 989;
        test_data[600] = 33'd6516032812;
        test_addr[601] = 990;
        test_data[601] = 33'd3379643487;
        test_addr[602] = 991;
        test_data[602] = 33'd6713643093;
        test_addr[603] = 992;
        test_data[603] = 33'd964179193;
        test_addr[604] = 993;
        test_data[604] = 33'd1857244546;
        test_addr[605] = 994;
        test_data[605] = 33'd7028511373;
        test_addr[606] = 995;
        test_data[606] = 33'd8040956289;
        test_addr[607] = 230;
        test_data[607] = 33'd2673908551;
        test_addr[608] = 231;
        test_data[608] = 33'd6051871487;
        test_addr[609] = 559;
        test_data[609] = 33'd839457297;
        test_addr[610] = 560;
        test_data[610] = 33'd2959208024;
        test_addr[611] = 561;
        test_data[611] = 33'd8173870982;
        test_addr[612] = 562;
        test_data[612] = 33'd1942238216;
        test_addr[613] = 563;
        test_data[613] = 33'd3656355596;
        test_addr[614] = 564;
        test_data[614] = 33'd1073823995;
        test_addr[615] = 565;
        test_data[615] = 33'd1483039500;
        test_addr[616] = 566;
        test_data[616] = 33'd3645197110;
        test_addr[617] = 232;
        test_data[617] = 33'd3657253458;
        test_addr[618] = 233;
        test_data[618] = 33'd5732469119;
        test_addr[619] = 234;
        test_data[619] = 33'd2569948806;
        test_addr[620] = 235;
        test_data[620] = 33'd2173127971;
        test_addr[621] = 236;
        test_data[621] = 33'd4837973217;
        test_addr[622] = 237;
        test_data[622] = 33'd2163671273;
        test_addr[623] = 238;
        test_data[623] = 33'd1309914105;
        test_addr[624] = 239;
        test_data[624] = 33'd5042423955;
        test_addr[625] = 240;
        test_data[625] = 33'd5859263288;
        test_addr[626] = 241;
        test_data[626] = 33'd738113948;
        test_addr[627] = 242;
        test_data[627] = 33'd5916344848;
        test_addr[628] = 243;
        test_data[628] = 33'd4757651253;
        test_addr[629] = 244;
        test_data[629] = 33'd3986444448;
        test_addr[630] = 245;
        test_data[630] = 33'd3509345496;
        test_addr[631] = 246;
        test_data[631] = 33'd2440705799;
        test_addr[632] = 247;
        test_data[632] = 33'd6497620364;
        test_addr[633] = 248;
        test_data[633] = 33'd5937542180;
        test_addr[634] = 249;
        test_data[634] = 33'd4121500431;
        test_addr[635] = 793;
        test_data[635] = 33'd1843129498;
        test_addr[636] = 794;
        test_data[636] = 33'd6205876210;
        test_addr[637] = 795;
        test_data[637] = 33'd1540072738;
        test_addr[638] = 796;
        test_data[638] = 33'd1292528924;
        test_addr[639] = 797;
        test_data[639] = 33'd5052889842;
        test_addr[640] = 798;
        test_data[640] = 33'd2831706730;
        test_addr[641] = 799;
        test_data[641] = 33'd1361996462;
        test_addr[642] = 800;
        test_data[642] = 33'd2684303926;
        test_addr[643] = 801;
        test_data[643] = 33'd2873799072;
        test_addr[644] = 802;
        test_data[644] = 33'd3491622919;
        test_addr[645] = 803;
        test_data[645] = 33'd3660731959;
        test_addr[646] = 804;
        test_data[646] = 33'd5284796402;
        test_addr[647] = 805;
        test_data[647] = 33'd341095953;
        test_addr[648] = 806;
        test_data[648] = 33'd3109763568;
        test_addr[649] = 807;
        test_data[649] = 33'd619472320;
        test_addr[650] = 808;
        test_data[650] = 33'd3811340329;
        test_addr[651] = 809;
        test_data[651] = 33'd3174497928;
        test_addr[652] = 810;
        test_data[652] = 33'd848075204;
        test_addr[653] = 811;
        test_data[653] = 33'd1022680166;
        test_addr[654] = 812;
        test_data[654] = 33'd732597252;
        test_addr[655] = 813;
        test_data[655] = 33'd2469749640;
        test_addr[656] = 814;
        test_data[656] = 33'd3911919694;
        test_addr[657] = 815;
        test_data[657] = 33'd4204391240;
        test_addr[658] = 816;
        test_data[658] = 33'd3714792815;
        test_addr[659] = 817;
        test_data[659] = 33'd3647515413;
        test_addr[660] = 818;
        test_data[660] = 33'd3263948359;
        test_addr[661] = 819;
        test_data[661] = 33'd2910897927;
        test_addr[662] = 820;
        test_data[662] = 33'd2587666766;
        test_addr[663] = 821;
        test_data[663] = 33'd3918583867;
        test_addr[664] = 822;
        test_data[664] = 33'd4808168146;
        test_addr[665] = 823;
        test_data[665] = 33'd3228310104;
        test_addr[666] = 824;
        test_data[666] = 33'd7519192697;
        test_addr[667] = 825;
        test_data[667] = 33'd3901277367;
        test_addr[668] = 826;
        test_data[668] = 33'd4876601476;
        test_addr[669] = 827;
        test_data[669] = 33'd1733846292;
        test_addr[670] = 828;
        test_data[670] = 33'd5314330040;
        test_addr[671] = 829;
        test_data[671] = 33'd1668879510;
        test_addr[672] = 830;
        test_data[672] = 33'd3958563769;
        test_addr[673] = 831;
        test_data[673] = 33'd1616713383;
        test_addr[674] = 832;
        test_data[674] = 33'd2891161115;
        test_addr[675] = 833;
        test_data[675] = 33'd1222734269;
        test_addr[676] = 834;
        test_data[676] = 33'd3031697508;
        test_addr[677] = 835;
        test_data[677] = 33'd6281450841;
        test_addr[678] = 836;
        test_data[678] = 33'd579485165;
        test_addr[679] = 837;
        test_data[679] = 33'd2561173077;
        test_addr[680] = 838;
        test_data[680] = 33'd2449081523;
        test_addr[681] = 839;
        test_data[681] = 33'd2174987116;
        test_addr[682] = 840;
        test_data[682] = 33'd7068440181;
        test_addr[683] = 841;
        test_data[683] = 33'd846659615;
        test_addr[684] = 842;
        test_data[684] = 33'd3536331538;
        test_addr[685] = 843;
        test_data[685] = 33'd1817785861;
        test_addr[686] = 844;
        test_data[686] = 33'd5851890036;
        test_addr[687] = 845;
        test_data[687] = 33'd7985853697;
        test_addr[688] = 846;
        test_data[688] = 33'd3605947957;
        test_addr[689] = 250;
        test_data[689] = 33'd6875169213;
        test_addr[690] = 251;
        test_data[690] = 33'd6122596006;
        test_addr[691] = 252;
        test_data[691] = 33'd6834434726;
        test_addr[692] = 253;
        test_data[692] = 33'd1046892784;
        test_addr[693] = 254;
        test_data[693] = 33'd893686890;
        test_addr[694] = 255;
        test_data[694] = 33'd738701221;
        test_addr[695] = 256;
        test_data[695] = 33'd6133002960;
        test_addr[696] = 257;
        test_data[696] = 33'd7361823853;
        test_addr[697] = 258;
        test_data[697] = 33'd5263159303;
        test_addr[698] = 465;
        test_data[698] = 33'd5371483420;
        test_addr[699] = 466;
        test_data[699] = 33'd3459645207;
        test_addr[700] = 467;
        test_data[700] = 33'd2537057546;
        test_addr[701] = 259;
        test_data[701] = 33'd3199409289;
        test_addr[702] = 260;
        test_data[702] = 33'd3784376997;
        test_addr[703] = 261;
        test_data[703] = 33'd3435254937;
        test_addr[704] = 262;
        test_data[704] = 33'd6258359478;
        test_addr[705] = 263;
        test_data[705] = 33'd1168259603;
        test_addr[706] = 264;
        test_data[706] = 33'd3017312274;
        test_addr[707] = 265;
        test_data[707] = 33'd4232753553;
        test_addr[708] = 266;
        test_data[708] = 33'd7967533778;
        test_addr[709] = 267;
        test_data[709] = 33'd6961747180;
        test_addr[710] = 268;
        test_data[710] = 33'd5173952642;
        test_addr[711] = 596;
        test_data[711] = 33'd8189195198;
        test_addr[712] = 597;
        test_data[712] = 33'd6509352106;
        test_addr[713] = 598;
        test_data[713] = 33'd133191090;
        test_addr[714] = 599;
        test_data[714] = 33'd7405506739;
        test_addr[715] = 600;
        test_data[715] = 33'd6379589289;
        test_addr[716] = 601;
        test_data[716] = 33'd1528966083;
        test_addr[717] = 602;
        test_data[717] = 33'd2985258556;
        test_addr[718] = 603;
        test_data[718] = 33'd1521945037;
        test_addr[719] = 604;
        test_data[719] = 33'd2635934467;
        test_addr[720] = 605;
        test_data[720] = 33'd6926084846;
        test_addr[721] = 606;
        test_data[721] = 33'd4613034254;
        test_addr[722] = 607;
        test_data[722] = 33'd3129915412;
        test_addr[723] = 608;
        test_data[723] = 33'd8509326600;
        test_addr[724] = 609;
        test_data[724] = 33'd2651952637;
        test_addr[725] = 269;
        test_data[725] = 33'd8033679110;
        test_addr[726] = 270;
        test_data[726] = 33'd5297123590;
        test_addr[727] = 271;
        test_data[727] = 33'd5309030378;
        test_addr[728] = 272;
        test_data[728] = 33'd8198558678;
        test_addr[729] = 273;
        test_data[729] = 33'd2852287615;
        test_addr[730] = 274;
        test_data[730] = 33'd3297475855;
        test_addr[731] = 275;
        test_data[731] = 33'd5997416981;
        test_addr[732] = 276;
        test_data[732] = 33'd151084863;
        test_addr[733] = 277;
        test_data[733] = 33'd1313409944;
        test_addr[734] = 278;
        test_data[734] = 33'd3951155712;
        test_addr[735] = 279;
        test_data[735] = 33'd2152272633;
        test_addr[736] = 280;
        test_data[736] = 33'd1318904363;
        test_addr[737] = 281;
        test_data[737] = 33'd1519219586;
        test_addr[738] = 282;
        test_data[738] = 33'd443030348;
        test_addr[739] = 283;
        test_data[739] = 33'd1573656911;
        test_addr[740] = 284;
        test_data[740] = 33'd8005567672;
        test_addr[741] = 285;
        test_data[741] = 33'd4078885917;
        test_addr[742] = 286;
        test_data[742] = 33'd7025539037;
        test_addr[743] = 287;
        test_data[743] = 33'd1630502931;
        test_addr[744] = 288;
        test_data[744] = 33'd5065089680;
        test_addr[745] = 289;
        test_data[745] = 33'd4555121833;
        test_addr[746] = 290;
        test_data[746] = 33'd7790227563;
        test_addr[747] = 711;
        test_data[747] = 33'd1104666845;
        test_addr[748] = 291;
        test_data[748] = 33'd4964893893;
        test_addr[749] = 292;
        test_data[749] = 33'd6645316564;
        test_addr[750] = 459;
        test_data[750] = 33'd826235681;
        test_addr[751] = 460;
        test_data[751] = 33'd3390313948;
        test_addr[752] = 461;
        test_data[752] = 33'd5875677308;
        test_addr[753] = 462;
        test_data[753] = 33'd3770112161;
        test_addr[754] = 463;
        test_data[754] = 33'd2623477901;
        test_addr[755] = 464;
        test_data[755] = 33'd3147145687;
        test_addr[756] = 465;
        test_data[756] = 33'd1076516124;
        test_addr[757] = 466;
        test_data[757] = 33'd3459645207;
        test_addr[758] = 467;
        test_data[758] = 33'd4945083915;
        test_addr[759] = 468;
        test_data[759] = 33'd3992930714;
        test_addr[760] = 469;
        test_data[760] = 33'd1664670904;
        test_addr[761] = 470;
        test_data[761] = 33'd7905297725;
        test_addr[762] = 471;
        test_data[762] = 33'd432895216;
        test_addr[763] = 472;
        test_data[763] = 33'd8102845968;
        test_addr[764] = 473;
        test_data[764] = 33'd1293966191;
        test_addr[765] = 474;
        test_data[765] = 33'd3708729244;
        test_addr[766] = 293;
        test_data[766] = 33'd880389596;
        test_addr[767] = 294;
        test_data[767] = 33'd6335875285;
        test_addr[768] = 295;
        test_data[768] = 33'd1453477040;
        test_addr[769] = 296;
        test_data[769] = 33'd72603561;
        test_addr[770] = 297;
        test_data[770] = 33'd5445169435;
        test_addr[771] = 298;
        test_data[771] = 33'd189733476;
        test_addr[772] = 299;
        test_data[772] = 33'd1004966428;
        test_addr[773] = 300;
        test_data[773] = 33'd1786211448;
        test_addr[774] = 301;
        test_data[774] = 33'd2613515428;
        test_addr[775] = 302;
        test_data[775] = 33'd3250392161;
        test_addr[776] = 303;
        test_data[776] = 33'd4095352313;
        test_addr[777] = 304;
        test_data[777] = 33'd3750445638;
        test_addr[778] = 99;
        test_data[778] = 33'd1718939551;
        test_addr[779] = 100;
        test_data[779] = 33'd3845605637;
        test_addr[780] = 101;
        test_data[780] = 33'd669798772;
        test_addr[781] = 102;
        test_data[781] = 33'd746597445;
        test_addr[782] = 103;
        test_data[782] = 33'd7537100195;
        test_addr[783] = 104;
        test_data[783] = 33'd5781362120;
        test_addr[784] = 105;
        test_data[784] = 33'd1511183284;
        test_addr[785] = 106;
        test_data[785] = 33'd8462053692;
        test_addr[786] = 107;
        test_data[786] = 33'd4002934247;
        test_addr[787] = 108;
        test_data[787] = 33'd1129779635;
        test_addr[788] = 109;
        test_data[788] = 33'd1300879613;
        test_addr[789] = 110;
        test_data[789] = 33'd1563193765;
        test_addr[790] = 305;
        test_data[790] = 33'd4667689711;
        test_addr[791] = 306;
        test_data[791] = 33'd7208946196;
        test_addr[792] = 307;
        test_data[792] = 33'd4030103948;
        test_addr[793] = 788;
        test_data[793] = 33'd3817033739;
        test_addr[794] = 789;
        test_data[794] = 33'd484067223;
        test_addr[795] = 790;
        test_data[795] = 33'd6222326350;
        test_addr[796] = 791;
        test_data[796] = 33'd505251469;
        test_addr[797] = 792;
        test_data[797] = 33'd3388575783;
        test_addr[798] = 793;
        test_data[798] = 33'd5308012460;
        test_addr[799] = 794;
        test_data[799] = 33'd1910908914;
        test_addr[800] = 795;
        test_data[800] = 33'd7040084613;
        test_addr[801] = 796;
        test_data[801] = 33'd7540882691;
        test_addr[802] = 797;
        test_data[802] = 33'd757922546;
        test_addr[803] = 798;
        test_data[803] = 33'd2831706730;
        test_addr[804] = 799;
        test_data[804] = 33'd6410147368;
        test_addr[805] = 800;
        test_data[805] = 33'd2684303926;
        test_addr[806] = 801;
        test_data[806] = 33'd2873799072;
        test_addr[807] = 802;
        test_data[807] = 33'd6216999222;
        test_addr[808] = 803;
        test_data[808] = 33'd3660731959;
        test_addr[809] = 804;
        test_data[809] = 33'd989829106;
        test_addr[810] = 805;
        test_data[810] = 33'd341095953;
        test_addr[811] = 806;
        test_data[811] = 33'd3109763568;
        test_addr[812] = 807;
        test_data[812] = 33'd619472320;
        test_addr[813] = 808;
        test_data[813] = 33'd3811340329;
        test_addr[814] = 809;
        test_data[814] = 33'd3174497928;
        test_addr[815] = 810;
        test_data[815] = 33'd848075204;
        test_addr[816] = 811;
        test_data[816] = 33'd1022680166;
        test_addr[817] = 812;
        test_data[817] = 33'd732597252;
        test_addr[818] = 813;
        test_data[818] = 33'd5534507367;
        test_addr[819] = 814;
        test_data[819] = 33'd7387739195;
        test_addr[820] = 815;
        test_data[820] = 33'd4204391240;
        test_addr[821] = 816;
        test_data[821] = 33'd5610362942;
        test_addr[822] = 817;
        test_data[822] = 33'd3647515413;
        test_addr[823] = 818;
        test_data[823] = 33'd8172854227;
        test_addr[824] = 819;
        test_data[824] = 33'd2910897927;
        test_addr[825] = 820;
        test_data[825] = 33'd8080541412;
        test_addr[826] = 821;
        test_data[826] = 33'd3918583867;
        test_addr[827] = 822;
        test_data[827] = 33'd4422411857;
        test_addr[828] = 823;
        test_data[828] = 33'd5638962959;
        test_addr[829] = 824;
        test_data[829] = 33'd3224225401;
        test_addr[830] = 825;
        test_data[830] = 33'd6900270226;
        test_addr[831] = 826;
        test_data[831] = 33'd581634180;
        test_addr[832] = 827;
        test_data[832] = 33'd6746701763;
        test_addr[833] = 308;
        test_data[833] = 33'd2797128928;
        test_addr[834] = 309;
        test_data[834] = 33'd1328657515;
        test_addr[835] = 310;
        test_data[835] = 33'd5891877079;
        test_addr[836] = 311;
        test_data[836] = 33'd3422864683;
        test_addr[837] = 312;
        test_data[837] = 33'd2136184510;
        test_addr[838] = 313;
        test_data[838] = 33'd3975800125;
        test_addr[839] = 314;
        test_data[839] = 33'd1771827745;
        test_addr[840] = 315;
        test_data[840] = 33'd5327575798;
        test_addr[841] = 316;
        test_data[841] = 33'd7256802397;
        test_addr[842] = 317;
        test_data[842] = 33'd613544344;
        test_addr[843] = 318;
        test_data[843] = 33'd5665388369;
        test_addr[844] = 319;
        test_data[844] = 33'd180363106;
        test_addr[845] = 320;
        test_data[845] = 33'd4010594226;
        test_addr[846] = 321;
        test_data[846] = 33'd6004763230;
        test_addr[847] = 322;
        test_data[847] = 33'd6545890039;
        test_addr[848] = 445;
        test_data[848] = 33'd1931819170;
        test_addr[849] = 446;
        test_data[849] = 33'd6312976080;
        test_addr[850] = 447;
        test_data[850] = 33'd1470049012;
        test_addr[851] = 448;
        test_data[851] = 33'd3836817188;
        test_addr[852] = 449;
        test_data[852] = 33'd4852820264;
        test_addr[853] = 450;
        test_data[853] = 33'd6066066264;
        test_addr[854] = 451;
        test_data[854] = 33'd6870590988;
        test_addr[855] = 452;
        test_data[855] = 33'd5644180599;
        test_addr[856] = 453;
        test_data[856] = 33'd3913516686;
        test_addr[857] = 454;
        test_data[857] = 33'd3918291114;
        test_addr[858] = 455;
        test_data[858] = 33'd5690463324;
        test_addr[859] = 456;
        test_data[859] = 33'd2655493248;
        test_addr[860] = 457;
        test_data[860] = 33'd2493953492;
        test_addr[861] = 323;
        test_data[861] = 33'd5994367764;
        test_addr[862] = 324;
        test_data[862] = 33'd4124680673;
        test_addr[863] = 325;
        test_data[863] = 33'd1292476535;
        test_addr[864] = 326;
        test_data[864] = 33'd3211040190;
        test_addr[865] = 327;
        test_data[865] = 33'd4021375997;
        test_addr[866] = 328;
        test_data[866] = 33'd7495049943;
        test_addr[867] = 329;
        test_data[867] = 33'd508970632;
        test_addr[868] = 330;
        test_data[868] = 33'd2871069657;
        test_addr[869] = 331;
        test_data[869] = 33'd3021584846;
        test_addr[870] = 332;
        test_data[870] = 33'd3802541065;
        test_addr[871] = 333;
        test_data[871] = 33'd3777587601;
        test_addr[872] = 334;
        test_data[872] = 33'd2560750633;
        test_addr[873] = 335;
        test_data[873] = 33'd3132902255;
        test_addr[874] = 336;
        test_data[874] = 33'd535597245;
        test_addr[875] = 337;
        test_data[875] = 33'd2803068549;
        test_addr[876] = 338;
        test_data[876] = 33'd1957293410;
        test_addr[877] = 517;
        test_data[877] = 33'd2393872258;
        test_addr[878] = 518;
        test_data[878] = 33'd5186968668;
        test_addr[879] = 519;
        test_data[879] = 33'd705002716;
        test_addr[880] = 520;
        test_data[880] = 33'd6485875875;
        test_addr[881] = 339;
        test_data[881] = 33'd8222322182;
        test_addr[882] = 340;
        test_data[882] = 33'd5375770055;
        test_addr[883] = 341;
        test_data[883] = 33'd3105826626;
        test_addr[884] = 342;
        test_data[884] = 33'd4307939510;
        test_addr[885] = 343;
        test_data[885] = 33'd3938949624;
        test_addr[886] = 344;
        test_data[886] = 33'd7082501256;
        test_addr[887] = 345;
        test_data[887] = 33'd4504856431;
        test_addr[888] = 346;
        test_data[888] = 33'd337408017;
        test_addr[889] = 347;
        test_data[889] = 33'd8392927338;
        test_addr[890] = 295;
        test_data[890] = 33'd7377711989;
        test_addr[891] = 296;
        test_data[891] = 33'd4419790671;
        test_addr[892] = 297;
        test_data[892] = 33'd5861503044;
        test_addr[893] = 298;
        test_data[893] = 33'd4721299615;
        test_addr[894] = 299;
        test_data[894] = 33'd1004966428;
        test_addr[895] = 300;
        test_data[895] = 33'd1786211448;
        test_addr[896] = 301;
        test_data[896] = 33'd4473091386;
        test_addr[897] = 302;
        test_data[897] = 33'd3250392161;
        test_addr[898] = 303;
        test_data[898] = 33'd7812133483;
        test_addr[899] = 304;
        test_data[899] = 33'd3750445638;
        test_addr[900] = 305;
        test_data[900] = 33'd6564069632;
        test_addr[901] = 306;
        test_data[901] = 33'd2913978900;
        test_addr[902] = 307;
        test_data[902] = 33'd4030103948;
        test_addr[903] = 308;
        test_data[903] = 33'd8544923012;
        test_addr[904] = 348;
        test_data[904] = 33'd3314453200;
        test_addr[905] = 349;
        test_data[905] = 33'd2590479583;
        test_addr[906] = 350;
        test_data[906] = 33'd5638433950;
        test_addr[907] = 351;
        test_data[907] = 33'd7128748049;
        test_addr[908] = 352;
        test_data[908] = 33'd5693896151;
        test_addr[909] = 635;
        test_data[909] = 33'd1607332002;
        test_addr[910] = 636;
        test_data[910] = 33'd2445663499;
        test_addr[911] = 637;
        test_data[911] = 33'd5300719877;
        test_addr[912] = 638;
        test_data[912] = 33'd4136659456;
        test_addr[913] = 639;
        test_data[913] = 33'd86901798;
        test_addr[914] = 640;
        test_data[914] = 33'd3316842311;
        test_addr[915] = 353;
        test_data[915] = 33'd4764615865;
        test_addr[916] = 354;
        test_data[916] = 33'd369923590;
        test_addr[917] = 355;
        test_data[917] = 33'd2603783369;
        test_addr[918] = 356;
        test_data[918] = 33'd5481395913;
        test_addr[919] = 357;
        test_data[919] = 33'd6146773141;
        test_addr[920] = 358;
        test_data[920] = 33'd3479819972;
        test_addr[921] = 359;
        test_data[921] = 33'd309287193;
        test_addr[922] = 360;
        test_data[922] = 33'd5066590507;
        test_addr[923] = 361;
        test_data[923] = 33'd2280030852;
        test_addr[924] = 362;
        test_data[924] = 33'd7046558305;
        test_addr[925] = 363;
        test_data[925] = 33'd3362159751;
        test_addr[926] = 364;
        test_data[926] = 33'd4091092656;
        test_addr[927] = 481;
        test_data[927] = 33'd3104519648;
        test_addr[928] = 482;
        test_data[928] = 33'd5236845891;
        test_addr[929] = 483;
        test_data[929] = 33'd7159034488;
        test_addr[930] = 484;
        test_data[930] = 33'd8401752809;
        test_addr[931] = 485;
        test_data[931] = 33'd3869014208;
        test_addr[932] = 486;
        test_data[932] = 33'd1136344694;
        test_addr[933] = 487;
        test_data[933] = 33'd5613416595;
        test_addr[934] = 488;
        test_data[934] = 33'd7197136116;
        test_addr[935] = 489;
        test_data[935] = 33'd7980949838;
        test_addr[936] = 490;
        test_data[936] = 33'd3475954419;
        test_addr[937] = 491;
        test_data[937] = 33'd2109522773;
        test_addr[938] = 492;
        test_data[938] = 33'd5906892491;
        test_addr[939] = 493;
        test_data[939] = 33'd8252411919;
        test_addr[940] = 494;
        test_data[940] = 33'd297707220;
        test_addr[941] = 495;
        test_data[941] = 33'd759490144;
        test_addr[942] = 496;
        test_data[942] = 33'd7761793546;
        test_addr[943] = 497;
        test_data[943] = 33'd1711199328;
        test_addr[944] = 498;
        test_data[944] = 33'd3738045385;
        test_addr[945] = 499;
        test_data[945] = 33'd4818359627;
        test_addr[946] = 500;
        test_data[946] = 33'd5287485299;
        test_addr[947] = 365;
        test_data[947] = 33'd7452163958;
        test_addr[948] = 366;
        test_data[948] = 33'd2904869292;
        test_addr[949] = 367;
        test_data[949] = 33'd5117369249;
        test_addr[950] = 368;
        test_data[950] = 33'd1594529834;
        test_addr[951] = 369;
        test_data[951] = 33'd1912926533;
        test_addr[952] = 370;
        test_data[952] = 33'd7510477758;
        test_addr[953] = 371;
        test_data[953] = 33'd1688419579;
        test_addr[954] = 372;
        test_data[954] = 33'd3823632809;
        test_addr[955] = 373;
        test_data[955] = 33'd3237219661;
        test_addr[956] = 374;
        test_data[956] = 33'd149363693;
        test_addr[957] = 375;
        test_data[957] = 33'd2093158352;
        test_addr[958] = 376;
        test_data[958] = 33'd736569085;
        test_addr[959] = 377;
        test_data[959] = 33'd1111968953;
        test_addr[960] = 378;
        test_data[960] = 33'd4089108044;
        test_addr[961] = 379;
        test_data[961] = 33'd2445988135;
        test_addr[962] = 380;
        test_data[962] = 33'd2614266083;
        test_addr[963] = 155;
        test_data[963] = 33'd1633875019;
        test_addr[964] = 156;
        test_data[964] = 33'd997076171;
        test_addr[965] = 157;
        test_data[965] = 33'd98365346;
        test_addr[966] = 158;
        test_data[966] = 33'd2430407245;
        test_addr[967] = 381;
        test_data[967] = 33'd3380814185;
        test_addr[968] = 382;
        test_data[968] = 33'd7289648699;
        test_addr[969] = 278;
        test_data[969] = 33'd3951155712;
        test_addr[970] = 279;
        test_data[970] = 33'd2152272633;
        test_addr[971] = 280;
        test_data[971] = 33'd4448652159;
        test_addr[972] = 383;
        test_data[972] = 33'd4756040729;
        test_addr[973] = 370;
        test_data[973] = 33'd3215510462;
        test_addr[974] = 371;
        test_data[974] = 33'd5391837300;
        test_addr[975] = 372;
        test_data[975] = 33'd3823632809;
        test_addr[976] = 373;
        test_data[976] = 33'd3237219661;
        test_addr[977] = 374;
        test_data[977] = 33'd149363693;
        test_addr[978] = 375;
        test_data[978] = 33'd2093158352;
        test_addr[979] = 376;
        test_data[979] = 33'd736569085;
        test_addr[980] = 377;
        test_data[980] = 33'd6851581659;
        test_addr[981] = 378;
        test_data[981] = 33'd4801095209;
        test_addr[982] = 379;
        test_data[982] = 33'd7583715475;
        test_addr[983] = 380;
        test_data[983] = 33'd2614266083;
        test_addr[984] = 381;
        test_data[984] = 33'd3380814185;
        test_addr[985] = 382;
        test_data[985] = 33'd2994681403;
        test_addr[986] = 384;
        test_data[986] = 33'd739005625;
        test_addr[987] = 385;
        test_data[987] = 33'd698224158;
        test_addr[988] = 386;
        test_data[988] = 33'd1877039969;
        test_addr[989] = 387;
        test_data[989] = 33'd140765230;
        test_addr[990] = 388;
        test_data[990] = 33'd8506587796;
        test_addr[991] = 389;
        test_data[991] = 33'd5425466698;
        test_addr[992] = 390;
        test_data[992] = 33'd2928158067;
        test_addr[993] = 391;
        test_data[993] = 33'd1779555079;
        test_addr[994] = 392;
        test_data[994] = 33'd10599762;
        test_addr[995] = 393;
        test_data[995] = 33'd1215078312;
        test_addr[996] = 394;
        test_data[996] = 33'd2899126994;
        test_addr[997] = 395;
        test_data[997] = 33'd4037953191;
        test_addr[998] = 396;
        test_data[998] = 33'd6516277583;
        test_addr[999] = 397;
        test_data[999] = 33'd3740595799;
        test_addr[1000] = 398;
        test_data[1000] = 33'd1885338136;
        test_addr[1001] = 399;
        test_data[1001] = 33'd798523023;
        test_addr[1002] = 400;
        test_data[1002] = 33'd12061985;
        test_addr[1003] = 401;
        test_data[1003] = 33'd1367308988;
        test_addr[1004] = 402;
        test_data[1004] = 33'd3328109157;
        test_addr[1005] = 403;
        test_data[1005] = 33'd1931821484;
        test_addr[1006] = 404;
        test_data[1006] = 33'd1720976526;
        test_addr[1007] = 405;
        test_data[1007] = 33'd7426646050;
        test_addr[1008] = 406;
        test_data[1008] = 33'd8399581589;
        test_addr[1009] = 407;
        test_data[1009] = 33'd3124378955;
        test_addr[1010] = 408;
        test_data[1010] = 33'd3784952382;
        test_addr[1011] = 409;
        test_data[1011] = 33'd829691805;
        test_addr[1012] = 410;
        test_data[1012] = 33'd1292454337;
        test_addr[1013] = 411;
        test_data[1013] = 33'd1053791089;
        test_addr[1014] = 1014;
        test_data[1014] = 33'd414447015;
        test_addr[1015] = 1015;
        test_data[1015] = 33'd4068782698;
        test_addr[1016] = 1016;
        test_data[1016] = 33'd6337169055;
        test_addr[1017] = 1017;
        test_data[1017] = 33'd3652225397;
        test_addr[1018] = 1018;
        test_data[1018] = 33'd2984861369;
        test_addr[1019] = 1019;
        test_data[1019] = 33'd5048241971;
        test_addr[1020] = 1020;
        test_data[1020] = 33'd4349403140;
        test_addr[1021] = 412;
        test_data[1021] = 33'd1038301027;
        test_addr[1022] = 413;
        test_data[1022] = 33'd2856665508;
        test_addr[1023] = 414;
        test_data[1023] = 33'd1136158832;
        test_addr[1024] = 415;
        test_data[1024] = 33'd268942874;
        test_addr[1025] = 416;
        test_data[1025] = 33'd2315947450;
        test_addr[1026] = 417;
        test_data[1026] = 33'd2168180925;
        test_addr[1027] = 418;
        test_data[1027] = 33'd7414094416;
        test_addr[1028] = 419;
        test_data[1028] = 33'd3511401386;
        test_addr[1029] = 420;
        test_data[1029] = 33'd2422752708;
        test_addr[1030] = 421;
        test_data[1030] = 33'd257964552;
        test_addr[1031] = 422;
        test_data[1031] = 33'd962672775;
        test_addr[1032] = 423;
        test_data[1032] = 33'd3728980285;
        test_addr[1033] = 424;
        test_data[1033] = 33'd4304180058;
        test_addr[1034] = 425;
        test_data[1034] = 33'd3494559305;
        test_addr[1035] = 426;
        test_data[1035] = 33'd3544872180;
        test_addr[1036] = 427;
        test_data[1036] = 33'd2561035456;
        test_addr[1037] = 428;
        test_data[1037] = 33'd3571198896;
        test_addr[1038] = 429;
        test_data[1038] = 33'd8545457988;
        test_addr[1039] = 430;
        test_data[1039] = 33'd5264612892;
        test_addr[1040] = 431;
        test_data[1040] = 33'd7084983338;
        test_addr[1041] = 432;
        test_data[1041] = 33'd3691339593;
        test_addr[1042] = 433;
        test_data[1042] = 33'd6294232260;
        test_addr[1043] = 234;
        test_data[1043] = 33'd2569948806;
        test_addr[1044] = 434;
        test_data[1044] = 33'd6306608993;
        test_addr[1045] = 435;
        test_data[1045] = 33'd6383886277;
        test_addr[1046] = 436;
        test_data[1046] = 33'd1804759271;
        test_addr[1047] = 437;
        test_data[1047] = 33'd446220078;
        test_addr[1048] = 438;
        test_data[1048] = 33'd943277004;
        test_addr[1049] = 1016;
        test_data[1049] = 33'd2042201759;
        test_addr[1050] = 1017;
        test_data[1050] = 33'd5086161904;
        test_addr[1051] = 1018;
        test_data[1051] = 33'd2984861369;
        test_addr[1052] = 1019;
        test_data[1052] = 33'd5477914456;
        test_addr[1053] = 1020;
        test_data[1053] = 33'd54435844;
        test_addr[1054] = 1021;
        test_data[1054] = 33'd229156893;
        test_addr[1055] = 1022;
        test_data[1055] = 33'd657762763;
        test_addr[1056] = 1023;
        test_data[1056] = 33'd2095860060;
        test_addr[1057] = 0;
        test_data[1057] = 33'd4892549877;
        test_addr[1058] = 1;
        test_data[1058] = 33'd7259384483;
        test_addr[1059] = 2;
        test_data[1059] = 33'd244488320;
        test_addr[1060] = 3;
        test_data[1060] = 33'd2009627834;
        test_addr[1061] = 4;
        test_data[1061] = 33'd1187404859;
        test_addr[1062] = 5;
        test_data[1062] = 33'd3400165079;
        test_addr[1063] = 439;
        test_data[1063] = 33'd1055579969;
        test_addr[1064] = 440;
        test_data[1064] = 33'd867078260;
        test_addr[1065] = 441;
        test_data[1065] = 33'd700898576;
        test_addr[1066] = 442;
        test_data[1066] = 33'd7186015262;
        test_addr[1067] = 443;
        test_data[1067] = 33'd1114978954;
        test_addr[1068] = 444;
        test_data[1068] = 33'd2972090766;
        test_addr[1069] = 445;
        test_data[1069] = 33'd6687068619;
        test_addr[1070] = 446;
        test_data[1070] = 33'd2018008784;
        test_addr[1071] = 447;
        test_data[1071] = 33'd1470049012;
        test_addr[1072] = 448;
        test_data[1072] = 33'd3836817188;
        test_addr[1073] = 449;
        test_data[1073] = 33'd557852968;
        test_addr[1074] = 935;
        test_data[1074] = 33'd2632191667;
        test_addr[1075] = 450;
        test_data[1075] = 33'd1771098968;
        test_addr[1076] = 451;
        test_data[1076] = 33'd6119337877;
        test_addr[1077] = 452;
        test_data[1077] = 33'd1349213303;
        test_addr[1078] = 453;
        test_data[1078] = 33'd3913516686;
        test_addr[1079] = 454;
        test_data[1079] = 33'd3918291114;
        test_addr[1080] = 455;
        test_data[1080] = 33'd1395496028;
        test_addr[1081] = 327;
        test_data[1081] = 33'd4021375997;
        test_addr[1082] = 328;
        test_data[1082] = 33'd3200082647;
        test_addr[1083] = 329;
        test_data[1083] = 33'd508970632;
        test_addr[1084] = 456;
        test_data[1084] = 33'd7781812664;
        test_addr[1085] = 457;
        test_data[1085] = 33'd2493953492;
        test_addr[1086] = 458;
        test_data[1086] = 33'd5128417806;
        test_addr[1087] = 459;
        test_data[1087] = 33'd826235681;
        test_addr[1088] = 460;
        test_data[1088] = 33'd3390313948;
        test_addr[1089] = 461;
        test_data[1089] = 33'd1580710012;
        test_addr[1090] = 462;
        test_data[1090] = 33'd3770112161;
        test_addr[1091] = 463;
        test_data[1091] = 33'd8305203690;
        test_addr[1092] = 464;
        test_data[1092] = 33'd3147145687;
        test_addr[1093] = 465;
        test_data[1093] = 33'd1076516124;
        test_addr[1094] = 466;
        test_data[1094] = 33'd3459645207;
        test_addr[1095] = 467;
        test_data[1095] = 33'd5558573046;
        test_addr[1096] = 468;
        test_data[1096] = 33'd3992930714;
        test_addr[1097] = 469;
        test_data[1097] = 33'd7981276458;
        test_addr[1098] = 470;
        test_data[1098] = 33'd5316270417;
        test_addr[1099] = 471;
        test_data[1099] = 33'd8400583615;
        test_addr[1100] = 472;
        test_data[1100] = 33'd3807878672;
        test_addr[1101] = 473;
        test_data[1101] = 33'd7946566176;
        test_addr[1102] = 474;
        test_data[1102] = 33'd5123201920;
        test_addr[1103] = 475;
        test_data[1103] = 33'd8291595347;
        test_addr[1104] = 476;
        test_data[1104] = 33'd3560019982;
        test_addr[1105] = 477;
        test_data[1105] = 33'd3221152013;
        test_addr[1106] = 478;
        test_data[1106] = 33'd1227762368;
        test_addr[1107] = 479;
        test_data[1107] = 33'd4566717228;
        test_addr[1108] = 480;
        test_data[1108] = 33'd5685594865;
        test_addr[1109] = 481;
        test_data[1109] = 33'd3104519648;
        test_addr[1110] = 482;
        test_data[1110] = 33'd941878595;
        test_addr[1111] = 483;
        test_data[1111] = 33'd7929480932;
        test_addr[1112] = 484;
        test_data[1112] = 33'd4106785513;
        test_addr[1113] = 275;
        test_data[1113] = 33'd1702449685;
        test_addr[1114] = 276;
        test_data[1114] = 33'd151084863;
        test_addr[1115] = 277;
        test_data[1115] = 33'd1313409944;
        test_addr[1116] = 278;
        test_data[1116] = 33'd3951155712;
        test_addr[1117] = 279;
        test_data[1117] = 33'd2152272633;
        test_addr[1118] = 280;
        test_data[1118] = 33'd7580793971;
        test_addr[1119] = 281;
        test_data[1119] = 33'd1519219586;
        test_addr[1120] = 282;
        test_data[1120] = 33'd443030348;
        test_addr[1121] = 283;
        test_data[1121] = 33'd1573656911;
        test_addr[1122] = 284;
        test_data[1122] = 33'd7337814103;
        test_addr[1123] = 285;
        test_data[1123] = 33'd4078885917;
        test_addr[1124] = 286;
        test_data[1124] = 33'd2730571741;
        test_addr[1125] = 287;
        test_data[1125] = 33'd6385286669;
        test_addr[1126] = 288;
        test_data[1126] = 33'd7495297979;
        test_addr[1127] = 289;
        test_data[1127] = 33'd260154537;
        test_addr[1128] = 290;
        test_data[1128] = 33'd7285540117;
        test_addr[1129] = 291;
        test_data[1129] = 33'd669926597;
        test_addr[1130] = 292;
        test_data[1130] = 33'd6258655764;
        test_addr[1131] = 293;
        test_data[1131] = 33'd880389596;
        test_addr[1132] = 294;
        test_data[1132] = 33'd8232181960;
        test_addr[1133] = 295;
        test_data[1133] = 33'd3082744693;
        test_addr[1134] = 296;
        test_data[1134] = 33'd124823375;
        test_addr[1135] = 297;
        test_data[1135] = 33'd7392717617;
        test_addr[1136] = 485;
        test_data[1136] = 33'd6581362066;
        test_addr[1137] = 486;
        test_data[1137] = 33'd1136344694;
        test_addr[1138] = 487;
        test_data[1138] = 33'd1318449299;
        test_addr[1139] = 488;
        test_data[1139] = 33'd2902168820;
        test_addr[1140] = 372;
        test_data[1140] = 33'd6222694922;
        test_addr[1141] = 373;
        test_data[1141] = 33'd7793441594;
        test_addr[1142] = 374;
        test_data[1142] = 33'd149363693;
        test_addr[1143] = 489;
        test_data[1143] = 33'd3685982542;
        test_addr[1144] = 490;
        test_data[1144] = 33'd3475954419;
        test_addr[1145] = 491;
        test_data[1145] = 33'd6324902197;
        test_addr[1146] = 1003;
        test_data[1146] = 33'd6561757125;
        test_addr[1147] = 1004;
        test_data[1147] = 33'd6394459761;
        test_addr[1148] = 492;
        test_data[1148] = 33'd4498979947;
        test_addr[1149] = 493;
        test_data[1149] = 33'd5303509650;
        test_addr[1150] = 494;
        test_data[1150] = 33'd297707220;
        test_addr[1151] = 495;
        test_data[1151] = 33'd759490144;
        test_addr[1152] = 496;
        test_data[1152] = 33'd4962270469;
        test_addr[1153] = 497;
        test_data[1153] = 33'd1711199328;
        test_addr[1154] = 498;
        test_data[1154] = 33'd3738045385;
        test_addr[1155] = 499;
        test_data[1155] = 33'd5411064374;
        test_addr[1156] = 500;
        test_data[1156] = 33'd992518003;
        test_addr[1157] = 501;
        test_data[1157] = 33'd1809835966;
        test_addr[1158] = 502;
        test_data[1158] = 33'd2391045745;
        test_addr[1159] = 503;
        test_data[1159] = 33'd6242444032;
        test_addr[1160] = 504;
        test_data[1160] = 33'd2260143172;
        test_addr[1161] = 505;
        test_data[1161] = 33'd6485866379;
        test_addr[1162] = 506;
        test_data[1162] = 33'd8583705751;
        test_addr[1163] = 507;
        test_data[1163] = 33'd724258612;
        test_addr[1164] = 508;
        test_data[1164] = 33'd5971279767;
        test_addr[1165] = 509;
        test_data[1165] = 33'd2006610656;
        test_addr[1166] = 283;
        test_data[1166] = 33'd4892309658;
        test_addr[1167] = 284;
        test_data[1167] = 33'd3042846807;
        test_addr[1168] = 285;
        test_data[1168] = 33'd4078885917;
        test_addr[1169] = 286;
        test_data[1169] = 33'd2730571741;
        test_addr[1170] = 287;
        test_data[1170] = 33'd8525954898;
        test_addr[1171] = 288;
        test_data[1171] = 33'd3200330683;
        test_addr[1172] = 289;
        test_data[1172] = 33'd6364967763;
        test_addr[1173] = 290;
        test_data[1173] = 33'd2990572821;
        test_addr[1174] = 291;
        test_data[1174] = 33'd669926597;
        test_addr[1175] = 292;
        test_data[1175] = 33'd1963688468;
        test_addr[1176] = 293;
        test_data[1176] = 33'd8383898841;
        test_addr[1177] = 294;
        test_data[1177] = 33'd3937214664;
        test_addr[1178] = 295;
        test_data[1178] = 33'd3082744693;
        test_addr[1179] = 296;
        test_data[1179] = 33'd124823375;
        test_addr[1180] = 297;
        test_data[1180] = 33'd7416247996;
        test_addr[1181] = 298;
        test_data[1181] = 33'd5882976869;
        test_addr[1182] = 299;
        test_data[1182] = 33'd1004966428;
        test_addr[1183] = 300;
        test_data[1183] = 33'd1786211448;
        test_addr[1184] = 301;
        test_data[1184] = 33'd178124090;
        test_addr[1185] = 302;
        test_data[1185] = 33'd3250392161;
        test_addr[1186] = 303;
        test_data[1186] = 33'd3517166187;
        test_addr[1187] = 304;
        test_data[1187] = 33'd6702934145;
        test_addr[1188] = 510;
        test_data[1188] = 33'd4129103904;
        test_addr[1189] = 511;
        test_data[1189] = 33'd1421325492;
        test_addr[1190] = 63;
        test_data[1190] = 33'd5724876230;
        test_addr[1191] = 64;
        test_data[1191] = 33'd3007627993;
        test_addr[1192] = 65;
        test_data[1192] = 33'd1673314307;
        test_addr[1193] = 66;
        test_data[1193] = 33'd4628717067;
        test_addr[1194] = 67;
        test_data[1194] = 33'd283800910;
        test_addr[1195] = 68;
        test_data[1195] = 33'd4896269692;
        test_addr[1196] = 69;
        test_data[1196] = 33'd7390980202;
        test_addr[1197] = 512;
        test_data[1197] = 33'd3788029954;
        test_addr[1198] = 513;
        test_data[1198] = 33'd4749903896;
        test_addr[1199] = 514;
        test_data[1199] = 33'd6321316260;
        test_addr[1200] = 515;
        test_data[1200] = 33'd2354318472;
        test_addr[1201] = 516;
        test_data[1201] = 33'd5004869087;
        test_addr[1202] = 517;
        test_data[1202] = 33'd2393872258;
        test_addr[1203] = 518;
        test_data[1203] = 33'd892001372;
        test_addr[1204] = 241;
        test_data[1204] = 33'd738113948;
        test_addr[1205] = 242;
        test_data[1205] = 33'd1621377552;
        test_addr[1206] = 243;
        test_data[1206] = 33'd7990848047;
        test_addr[1207] = 244;
        test_data[1207] = 33'd3986444448;
        test_addr[1208] = 245;
        test_data[1208] = 33'd7095363608;
        test_addr[1209] = 246;
        test_data[1209] = 33'd2440705799;
        test_addr[1210] = 247;
        test_data[1210] = 33'd5185530902;
        test_addr[1211] = 248;
        test_data[1211] = 33'd6630325174;
        test_addr[1212] = 249;
        test_data[1212] = 33'd5297805254;
        test_addr[1213] = 250;
        test_data[1213] = 33'd2580201917;
        test_addr[1214] = 251;
        test_data[1214] = 33'd1827628710;
        test_addr[1215] = 519;
        test_data[1215] = 33'd705002716;
        test_addr[1216] = 520;
        test_data[1216] = 33'd2190908579;
        test_addr[1217] = 521;
        test_data[1217] = 33'd1306264201;
        test_addr[1218] = 522;
        test_data[1218] = 33'd4806727829;
        test_addr[1219] = 523;
        test_data[1219] = 33'd1659053730;
        test_addr[1220] = 524;
        test_data[1220] = 33'd2535488802;
        test_addr[1221] = 525;
        test_data[1221] = 33'd6662522664;
        test_addr[1222] = 526;
        test_data[1222] = 33'd6813109563;
        test_addr[1223] = 527;
        test_data[1223] = 33'd3043177996;
        test_addr[1224] = 528;
        test_data[1224] = 33'd1208414750;
        test_addr[1225] = 529;
        test_data[1225] = 33'd1896802361;
        test_addr[1226] = 530;
        test_data[1226] = 33'd1192716121;
        test_addr[1227] = 531;
        test_data[1227] = 33'd4886776374;
        test_addr[1228] = 532;
        test_data[1228] = 33'd1329842884;
        test_addr[1229] = 533;
        test_data[1229] = 33'd4525555214;
        test_addr[1230] = 587;
        test_data[1230] = 33'd3912203569;
        test_addr[1231] = 588;
        test_data[1231] = 33'd2997617910;
        test_addr[1232] = 534;
        test_data[1232] = 33'd1623632665;
        test_addr[1233] = 535;
        test_data[1233] = 33'd5382576912;
        test_addr[1234] = 536;
        test_data[1234] = 33'd5896363318;
        test_addr[1235] = 537;
        test_data[1235] = 33'd6474987007;
        test_addr[1236] = 722;
        test_data[1236] = 33'd4264062206;
        test_addr[1237] = 723;
        test_data[1237] = 33'd2035228107;
        test_addr[1238] = 724;
        test_data[1238] = 33'd3488346519;
        test_addr[1239] = 725;
        test_data[1239] = 33'd4023969800;
        test_addr[1240] = 726;
        test_data[1240] = 33'd7358878438;
        test_addr[1241] = 727;
        test_data[1241] = 33'd2168181148;
        test_addr[1242] = 538;
        test_data[1242] = 33'd7503001257;
        test_addr[1243] = 539;
        test_data[1243] = 33'd6368462319;
        test_addr[1244] = 540;
        test_data[1244] = 33'd8026290638;
        test_addr[1245] = 541;
        test_data[1245] = 33'd1920105602;
        test_addr[1246] = 542;
        test_data[1246] = 33'd3693452330;
        test_addr[1247] = 543;
        test_data[1247] = 33'd1931463624;
        test_addr[1248] = 544;
        test_data[1248] = 33'd118999468;
        test_addr[1249] = 929;
        test_data[1249] = 33'd1467497009;
        test_addr[1250] = 545;
        test_data[1250] = 33'd1749290836;
        test_addr[1251] = 546;
        test_data[1251] = 33'd717909476;
        test_addr[1252] = 547;
        test_data[1252] = 33'd1656097789;
        test_addr[1253] = 548;
        test_data[1253] = 33'd3975122350;
        test_addr[1254] = 549;
        test_data[1254] = 33'd2127589844;
        test_addr[1255] = 550;
        test_data[1255] = 33'd3378215821;
        test_addr[1256] = 551;
        test_data[1256] = 33'd3550124624;
        test_addr[1257] = 552;
        test_data[1257] = 33'd1286678884;
        test_addr[1258] = 553;
        test_data[1258] = 33'd1687299562;
        test_addr[1259] = 554;
        test_data[1259] = 33'd5344546632;
        test_addr[1260] = 555;
        test_data[1260] = 33'd2248499919;
        test_addr[1261] = 556;
        test_data[1261] = 33'd2939472687;
        test_addr[1262] = 557;
        test_data[1262] = 33'd985122537;
        test_addr[1263] = 558;
        test_data[1263] = 33'd3808977718;
        test_addr[1264] = 559;
        test_data[1264] = 33'd839457297;
        test_addr[1265] = 427;
        test_data[1265] = 33'd5585562811;
        test_addr[1266] = 428;
        test_data[1266] = 33'd3571198896;
        test_addr[1267] = 429;
        test_data[1267] = 33'd4250490692;
        test_addr[1268] = 430;
        test_data[1268] = 33'd5238128759;
        test_addr[1269] = 431;
        test_data[1269] = 33'd2790016042;
        test_addr[1270] = 432;
        test_data[1270] = 33'd3691339593;
        test_addr[1271] = 433;
        test_data[1271] = 33'd1999264964;
        test_addr[1272] = 434;
        test_data[1272] = 33'd2011641697;
        test_addr[1273] = 435;
        test_data[1273] = 33'd2088918981;
        test_addr[1274] = 436;
        test_data[1274] = 33'd6946121856;
        test_addr[1275] = 560;
        test_data[1275] = 33'd5108702818;
        test_addr[1276] = 561;
        test_data[1276] = 33'd3878903686;
        test_addr[1277] = 562;
        test_data[1277] = 33'd1942238216;
        test_addr[1278] = 563;
        test_data[1278] = 33'd3656355596;
        test_addr[1279] = 564;
        test_data[1279] = 33'd4514783739;
        test_addr[1280] = 565;
        test_data[1280] = 33'd5437237978;
        test_addr[1281] = 566;
        test_data[1281] = 33'd7562921377;
        test_addr[1282] = 567;
        test_data[1282] = 33'd3156642332;
        test_addr[1283] = 568;
        test_data[1283] = 33'd148205842;
        test_addr[1284] = 569;
        test_data[1284] = 33'd4106722886;
        test_addr[1285] = 570;
        test_data[1285] = 33'd5046595994;
        test_addr[1286] = 540;
        test_data[1286] = 33'd7355299523;
        test_addr[1287] = 541;
        test_data[1287] = 33'd6137745499;
        test_addr[1288] = 542;
        test_data[1288] = 33'd3693452330;
        test_addr[1289] = 543;
        test_data[1289] = 33'd1931463624;
        test_addr[1290] = 544;
        test_data[1290] = 33'd118999468;
        test_addr[1291] = 545;
        test_data[1291] = 33'd7883706532;
        test_addr[1292] = 546;
        test_data[1292] = 33'd717909476;
        test_addr[1293] = 547;
        test_data[1293] = 33'd1656097789;
        test_addr[1294] = 548;
        test_data[1294] = 33'd3975122350;
        test_addr[1295] = 549;
        test_data[1295] = 33'd2127589844;
        test_addr[1296] = 550;
        test_data[1296] = 33'd3378215821;
        test_addr[1297] = 551;
        test_data[1297] = 33'd3550124624;
        test_addr[1298] = 552;
        test_data[1298] = 33'd5510165499;
        test_addr[1299] = 571;
        test_data[1299] = 33'd4031278286;
        test_addr[1300] = 572;
        test_data[1300] = 33'd7881349985;
        test_addr[1301] = 573;
        test_data[1301] = 33'd8087758049;
        test_addr[1302] = 574;
        test_data[1302] = 33'd5729214465;
        test_addr[1303] = 575;
        test_data[1303] = 33'd5776598225;
        test_addr[1304] = 576;
        test_data[1304] = 33'd7680048815;
        test_addr[1305] = 577;
        test_data[1305] = 33'd513421463;
        test_addr[1306] = 90;
        test_data[1306] = 33'd43380869;
        test_addr[1307] = 91;
        test_data[1307] = 33'd138001890;
        test_addr[1308] = 92;
        test_data[1308] = 33'd403469968;
        test_addr[1309] = 93;
        test_data[1309] = 33'd563973034;
        test_addr[1310] = 94;
        test_data[1310] = 33'd4213193887;
        test_addr[1311] = 95;
        test_data[1311] = 33'd610452162;
        test_addr[1312] = 96;
        test_data[1312] = 33'd8025479429;
        test_addr[1313] = 97;
        test_data[1313] = 33'd654962339;
        test_addr[1314] = 98;
        test_data[1314] = 33'd7084453552;
        test_addr[1315] = 99;
        test_data[1315] = 33'd1718939551;
        test_addr[1316] = 100;
        test_data[1316] = 33'd3845605637;
        test_addr[1317] = 578;
        test_data[1317] = 33'd2894820147;
        test_addr[1318] = 579;
        test_data[1318] = 33'd3224225652;
        test_addr[1319] = 909;
        test_data[1319] = 33'd6257557414;
        test_addr[1320] = 910;
        test_data[1320] = 33'd885454967;
        test_addr[1321] = 911;
        test_data[1321] = 33'd6234170121;
        test_addr[1322] = 912;
        test_data[1322] = 33'd5157601176;
        test_addr[1323] = 913;
        test_data[1323] = 33'd3108154670;
        test_addr[1324] = 580;
        test_data[1324] = 33'd1239202064;
        test_addr[1325] = 581;
        test_data[1325] = 33'd5744041671;
        test_addr[1326] = 582;
        test_data[1326] = 33'd8123131333;
        test_addr[1327] = 583;
        test_data[1327] = 33'd5263626996;
        test_addr[1328] = 584;
        test_data[1328] = 33'd7485726537;
        test_addr[1329] = 712;
        test_data[1329] = 33'd3993640537;
        test_addr[1330] = 713;
        test_data[1330] = 33'd3877347980;
        test_addr[1331] = 714;
        test_data[1331] = 33'd1793666688;
        test_addr[1332] = 715;
        test_data[1332] = 33'd701885885;
        test_addr[1333] = 716;
        test_data[1333] = 33'd2594539979;
        test_addr[1334] = 717;
        test_data[1334] = 33'd6921151969;
        test_addr[1335] = 718;
        test_data[1335] = 33'd5601089114;
        test_addr[1336] = 719;
        test_data[1336] = 33'd3591465327;
        test_addr[1337] = 720;
        test_data[1337] = 33'd2657030068;
        test_addr[1338] = 721;
        test_data[1338] = 33'd662721243;
        test_addr[1339] = 585;
        test_data[1339] = 33'd4604120204;
        test_addr[1340] = 586;
        test_data[1340] = 33'd3389351130;
        test_addr[1341] = 587;
        test_data[1341] = 33'd3912203569;
        test_addr[1342] = 588;
        test_data[1342] = 33'd2997617910;
        test_addr[1343] = 589;
        test_data[1343] = 33'd788551438;
        test_addr[1344] = 590;
        test_data[1344] = 33'd7444752537;
        test_addr[1345] = 591;
        test_data[1345] = 33'd8113771672;
        test_addr[1346] = 592;
        test_data[1346] = 33'd3656952568;
        test_addr[1347] = 593;
        test_data[1347] = 33'd8393691248;
        test_addr[1348] = 594;
        test_data[1348] = 33'd2232370504;
        test_addr[1349] = 595;
        test_data[1349] = 33'd7739820636;
        test_addr[1350] = 596;
        test_data[1350] = 33'd3894227902;
        test_addr[1351] = 597;
        test_data[1351] = 33'd2214384810;
        test_addr[1352] = 598;
        test_data[1352] = 33'd133191090;
        test_addr[1353] = 599;
        test_data[1353] = 33'd6516698752;
        test_addr[1354] = 600;
        test_data[1354] = 33'd2084621993;
        test_addr[1355] = 601;
        test_data[1355] = 33'd1528966083;
        test_addr[1356] = 602;
        test_data[1356] = 33'd2985258556;
        test_addr[1357] = 603;
        test_data[1357] = 33'd1521945037;
        test_addr[1358] = 815;
        test_data[1358] = 33'd5161584303;
        test_addr[1359] = 816;
        test_data[1359] = 33'd1315395646;
        test_addr[1360] = 817;
        test_data[1360] = 33'd5083886202;
        test_addr[1361] = 818;
        test_data[1361] = 33'd3877886931;
        test_addr[1362] = 819;
        test_data[1362] = 33'd2910897927;
        test_addr[1363] = 820;
        test_data[1363] = 33'd5890800863;
        test_addr[1364] = 821;
        test_data[1364] = 33'd8238873364;
        test_addr[1365] = 822;
        test_data[1365] = 33'd6817170750;
        test_addr[1366] = 823;
        test_data[1366] = 33'd1343995663;
        test_addr[1367] = 824;
        test_data[1367] = 33'd3224225401;
        test_addr[1368] = 825;
        test_data[1368] = 33'd2605302930;
        test_addr[1369] = 826;
        test_data[1369] = 33'd581634180;
        test_addr[1370] = 827;
        test_data[1370] = 33'd4460848584;
        test_addr[1371] = 828;
        test_data[1371] = 33'd1019362744;
        test_addr[1372] = 829;
        test_data[1372] = 33'd1668879510;
        test_addr[1373] = 830;
        test_data[1373] = 33'd3958563769;
        test_addr[1374] = 831;
        test_data[1374] = 33'd1616713383;
        test_addr[1375] = 832;
        test_data[1375] = 33'd2891161115;
        test_addr[1376] = 604;
        test_data[1376] = 33'd6838748680;
        test_addr[1377] = 605;
        test_data[1377] = 33'd2631117550;
        test_addr[1378] = 606;
        test_data[1378] = 33'd318066958;
        test_addr[1379] = 607;
        test_data[1379] = 33'd3129915412;
        test_addr[1380] = 608;
        test_data[1380] = 33'd5377095208;
        test_addr[1381] = 609;
        test_data[1381] = 33'd2651952637;
        test_addr[1382] = 610;
        test_data[1382] = 33'd2655954426;
        test_addr[1383] = 611;
        test_data[1383] = 33'd507597236;
        test_addr[1384] = 612;
        test_data[1384] = 33'd3082247360;
        test_addr[1385] = 613;
        test_data[1385] = 33'd8212782335;
        test_addr[1386] = 614;
        test_data[1386] = 33'd4733190884;
        test_addr[1387] = 615;
        test_data[1387] = 33'd3553517321;
        test_addr[1388] = 616;
        test_data[1388] = 33'd1763094828;
        test_addr[1389] = 617;
        test_data[1389] = 33'd8589635760;
        test_addr[1390] = 618;
        test_data[1390] = 33'd2989005313;
        test_addr[1391] = 619;
        test_data[1391] = 33'd2093912685;
        test_addr[1392] = 620;
        test_data[1392] = 33'd7564720650;
        test_addr[1393] = 621;
        test_data[1393] = 33'd7011379347;
        test_addr[1394] = 622;
        test_data[1394] = 33'd5687034626;
        test_addr[1395] = 623;
        test_data[1395] = 33'd2296683503;
        test_addr[1396] = 624;
        test_data[1396] = 33'd50566768;
        test_addr[1397] = 625;
        test_data[1397] = 33'd3238708872;
        test_addr[1398] = 626;
        test_data[1398] = 33'd489015939;
        test_addr[1399] = 627;
        test_data[1399] = 33'd4452856415;
        test_addr[1400] = 628;
        test_data[1400] = 33'd2298215631;
        test_addr[1401] = 629;
        test_data[1401] = 33'd4372517962;
        test_addr[1402] = 630;
        test_data[1402] = 33'd4424045716;
        test_addr[1403] = 631;
        test_data[1403] = 33'd793101746;
        test_addr[1404] = 632;
        test_data[1404] = 33'd6251595718;
        test_addr[1405] = 633;
        test_data[1405] = 33'd7874238597;
        test_addr[1406] = 634;
        test_data[1406] = 33'd2429702712;
        test_addr[1407] = 635;
        test_data[1407] = 33'd1607332002;
        test_addr[1408] = 636;
        test_data[1408] = 33'd6634986565;
        test_addr[1409] = 1006;
        test_data[1409] = 33'd2573864613;
        test_addr[1410] = 637;
        test_data[1410] = 33'd1005752581;
        test_addr[1411] = 638;
        test_data[1411] = 33'd4136659456;
        test_addr[1412] = 639;
        test_data[1412] = 33'd86901798;
        test_addr[1413] = 640;
        test_data[1413] = 33'd5760952593;
        test_addr[1414] = 641;
        test_data[1414] = 33'd3586386131;
        test_addr[1415] = 642;
        test_data[1415] = 33'd5057137962;
        test_addr[1416] = 643;
        test_data[1416] = 33'd1955210064;
        test_addr[1417] = 644;
        test_data[1417] = 33'd2998446653;
        test_addr[1418] = 645;
        test_data[1418] = 33'd1474811439;
        test_addr[1419] = 646;
        test_data[1419] = 33'd1560612810;
        test_addr[1420] = 647;
        test_data[1420] = 33'd6641201661;
        test_addr[1421] = 648;
        test_data[1421] = 33'd2360713956;
        test_addr[1422] = 649;
        test_data[1422] = 33'd3349786723;
        test_addr[1423] = 650;
        test_data[1423] = 33'd4203221935;
        test_addr[1424] = 651;
        test_data[1424] = 33'd3706032235;
        test_addr[1425] = 652;
        test_data[1425] = 33'd7875677124;
        test_addr[1426] = 653;
        test_data[1426] = 33'd923572889;
        test_addr[1427] = 654;
        test_data[1427] = 33'd3014930614;
        test_addr[1428] = 601;
        test_data[1428] = 33'd1528966083;
        test_addr[1429] = 655;
        test_data[1429] = 33'd88765548;
        test_addr[1430] = 656;
        test_data[1430] = 33'd2492457321;
        test_addr[1431] = 657;
        test_data[1431] = 33'd576451002;
        test_addr[1432] = 658;
        test_data[1432] = 33'd171564132;
        test_addr[1433] = 659;
        test_data[1433] = 33'd4136402978;
        test_addr[1434] = 660;
        test_data[1434] = 33'd2157180827;
        test_addr[1435] = 661;
        test_data[1435] = 33'd5699460116;
        test_addr[1436] = 662;
        test_data[1436] = 33'd4126887004;
        test_addr[1437] = 663;
        test_data[1437] = 33'd3355262986;
        test_addr[1438] = 664;
        test_data[1438] = 33'd6714045190;
        test_addr[1439] = 665;
        test_data[1439] = 33'd998667060;
        test_addr[1440] = 666;
        test_data[1440] = 33'd4045379889;
        test_addr[1441] = 667;
        test_data[1441] = 33'd1268036190;
        test_addr[1442] = 668;
        test_data[1442] = 33'd1574161429;
        test_addr[1443] = 669;
        test_data[1443] = 33'd3372123763;
        test_addr[1444] = 670;
        test_data[1444] = 33'd2901628700;
        test_addr[1445] = 671;
        test_data[1445] = 33'd7985015171;
        test_addr[1446] = 672;
        test_data[1446] = 33'd3355015249;
        test_addr[1447] = 673;
        test_data[1447] = 33'd7699201383;
        test_addr[1448] = 674;
        test_data[1448] = 33'd2390983344;
        test_addr[1449] = 675;
        test_data[1449] = 33'd2709261325;
        test_addr[1450] = 676;
        test_data[1450] = 33'd1104785019;
        test_addr[1451] = 677;
        test_data[1451] = 33'd5224835122;
        test_addr[1452] = 488;
        test_data[1452] = 33'd2902168820;
        test_addr[1453] = 678;
        test_data[1453] = 33'd5531318348;
        test_addr[1454] = 253;
        test_data[1454] = 33'd1046892784;
        test_addr[1455] = 679;
        test_data[1455] = 33'd7971388478;
        test_addr[1456] = 680;
        test_data[1456] = 33'd3119041072;
        test_addr[1457] = 919;
        test_data[1457] = 33'd2511923435;
        test_addr[1458] = 920;
        test_data[1458] = 33'd3915123610;
        test_addr[1459] = 921;
        test_data[1459] = 33'd3532290497;
        test_addr[1460] = 922;
        test_data[1460] = 33'd181860439;
        test_addr[1461] = 923;
        test_data[1461] = 33'd5699241361;
        test_addr[1462] = 924;
        test_data[1462] = 33'd5505796954;
        test_addr[1463] = 925;
        test_data[1463] = 33'd1313195782;
        test_addr[1464] = 926;
        test_data[1464] = 33'd7879200910;
        test_addr[1465] = 927;
        test_data[1465] = 33'd877988174;
        test_addr[1466] = 928;
        test_data[1466] = 33'd3715639018;
        test_addr[1467] = 681;
        test_data[1467] = 33'd5991029629;
        test_addr[1468] = 682;
        test_data[1468] = 33'd6512946141;
        test_addr[1469] = 683;
        test_data[1469] = 33'd3097106317;
        test_addr[1470] = 684;
        test_data[1470] = 33'd1377128895;
        test_addr[1471] = 111;
        test_data[1471] = 33'd59269632;
        test_addr[1472] = 685;
        test_data[1472] = 33'd992539895;
        test_addr[1473] = 686;
        test_data[1473] = 33'd626729407;
        test_addr[1474] = 687;
        test_data[1474] = 33'd2332656559;
        test_addr[1475] = 688;
        test_data[1475] = 33'd6255613051;
        test_addr[1476] = 689;
        test_data[1476] = 33'd7115495832;
        test_addr[1477] = 690;
        test_data[1477] = 33'd1799699601;
        test_addr[1478] = 691;
        test_data[1478] = 33'd8209452529;
        test_addr[1479] = 692;
        test_data[1479] = 33'd5302299721;
        test_addr[1480] = 693;
        test_data[1480] = 33'd1755618517;
        test_addr[1481] = 694;
        test_data[1481] = 33'd1783902209;
        test_addr[1482] = 807;
        test_data[1482] = 33'd619472320;
        test_addr[1483] = 808;
        test_data[1483] = 33'd3811340329;
        test_addr[1484] = 809;
        test_data[1484] = 33'd3174497928;
        test_addr[1485] = 810;
        test_data[1485] = 33'd848075204;
        test_addr[1486] = 811;
        test_data[1486] = 33'd1022680166;
        test_addr[1487] = 812;
        test_data[1487] = 33'd5309588295;
        test_addr[1488] = 695;
        test_data[1488] = 33'd4120276502;
        test_addr[1489] = 696;
        test_data[1489] = 33'd1053390424;
        test_addr[1490] = 697;
        test_data[1490] = 33'd6968123720;
        test_addr[1491] = 698;
        test_data[1491] = 33'd8195369717;
        test_addr[1492] = 699;
        test_data[1492] = 33'd2973118482;
        test_addr[1493] = 700;
        test_data[1493] = 33'd968388609;
        test_addr[1494] = 701;
        test_data[1494] = 33'd835744670;
        test_addr[1495] = 640;
        test_data[1495] = 33'd1465985297;
        test_addr[1496] = 641;
        test_data[1496] = 33'd3586386131;
        test_addr[1497] = 642;
        test_data[1497] = 33'd762170666;
        test_addr[1498] = 643;
        test_data[1498] = 33'd4523543743;
        test_addr[1499] = 644;
        test_data[1499] = 33'd7977968766;
        test_addr[1500] = 645;
        test_data[1500] = 33'd1474811439;
        test_addr[1501] = 646;
        test_data[1501] = 33'd1560612810;
        test_addr[1502] = 647;
        test_data[1502] = 33'd2346234365;
        test_addr[1503] = 648;
        test_data[1503] = 33'd7356458099;
        test_addr[1504] = 702;
        test_data[1504] = 33'd5859695857;
        test_addr[1505] = 703;
        test_data[1505] = 33'd1255659046;
        test_addr[1506] = 704;
        test_data[1506] = 33'd998116682;
        test_addr[1507] = 705;
        test_data[1507] = 33'd1911257944;
        test_addr[1508] = 706;
        test_data[1508] = 33'd3521378079;
        test_addr[1509] = 707;
        test_data[1509] = 33'd7336621843;
        test_addr[1510] = 708;
        test_data[1510] = 33'd3884518045;
        test_addr[1511] = 709;
        test_data[1511] = 33'd3130440955;
        test_addr[1512] = 710;
        test_data[1512] = 33'd3654683160;
        test_addr[1513] = 711;
        test_data[1513] = 33'd7362927195;
        test_addr[1514] = 712;
        test_data[1514] = 33'd3993640537;
        test_addr[1515] = 713;
        test_data[1515] = 33'd3877347980;
        test_addr[1516] = 88;
        test_data[1516] = 33'd4739025778;
        test_addr[1517] = 89;
        test_data[1517] = 33'd461104171;
        test_addr[1518] = 90;
        test_data[1518] = 33'd43380869;
        test_addr[1519] = 714;
        test_data[1519] = 33'd1793666688;
        test_addr[1520] = 715;
        test_data[1520] = 33'd701885885;
        test_addr[1521] = 716;
        test_data[1521] = 33'd2594539979;
        test_addr[1522] = 717;
        test_data[1522] = 33'd2626184673;
        test_addr[1523] = 718;
        test_data[1523] = 33'd1306121818;
        test_addr[1524] = 719;
        test_data[1524] = 33'd3591465327;
        test_addr[1525] = 720;
        test_data[1525] = 33'd2657030068;
        test_addr[1526] = 721;
        test_data[1526] = 33'd662721243;
        test_addr[1527] = 722;
        test_data[1527] = 33'd4264062206;
        test_addr[1528] = 723;
        test_data[1528] = 33'd2035228107;
        test_addr[1529] = 724;
        test_data[1529] = 33'd3488346519;
        test_addr[1530] = 725;
        test_data[1530] = 33'd4023969800;
        test_addr[1531] = 726;
        test_data[1531] = 33'd3063911142;
        test_addr[1532] = 727;
        test_data[1532] = 33'd8521940929;
        test_addr[1533] = 728;
        test_data[1533] = 33'd716320088;
        test_addr[1534] = 729;
        test_data[1534] = 33'd5259574815;
        test_addr[1535] = 730;
        test_data[1535] = 33'd3458672318;
        test_addr[1536] = 731;
        test_data[1536] = 33'd1618801135;
        test_addr[1537] = 732;
        test_data[1537] = 33'd5186905860;
        test_addr[1538] = 144;
        test_data[1538] = 33'd4076204621;
        test_addr[1539] = 733;
        test_data[1539] = 33'd844566830;
        test_addr[1540] = 734;
        test_data[1540] = 33'd1357887344;
        test_addr[1541] = 735;
        test_data[1541] = 33'd5792048832;
        test_addr[1542] = 992;
        test_data[1542] = 33'd964179193;
        test_addr[1543] = 993;
        test_data[1543] = 33'd5643540822;
        test_addr[1544] = 994;
        test_data[1544] = 33'd2733544077;
        test_addr[1545] = 995;
        test_data[1545] = 33'd3745988993;
        test_addr[1546] = 996;
        test_data[1546] = 33'd3922015050;
        test_addr[1547] = 997;
        test_data[1547] = 33'd1759334156;
        test_addr[1548] = 998;
        test_data[1548] = 33'd6122676213;
        test_addr[1549] = 999;
        test_data[1549] = 33'd6399314956;
        test_addr[1550] = 736;
        test_data[1550] = 33'd914072280;
        test_addr[1551] = 737;
        test_data[1551] = 33'd565879052;
        test_addr[1552] = 738;
        test_data[1552] = 33'd3739241179;
        test_addr[1553] = 739;
        test_data[1553] = 33'd6572005514;
        test_addr[1554] = 740;
        test_data[1554] = 33'd2567066062;
        test_addr[1555] = 741;
        test_data[1555] = 33'd2013379092;
        test_addr[1556] = 742;
        test_data[1556] = 33'd546339758;
        test_addr[1557] = 743;
        test_data[1557] = 33'd2720583043;
        test_addr[1558] = 744;
        test_data[1558] = 33'd4202166401;
        test_addr[1559] = 745;
        test_data[1559] = 33'd6533691328;
        test_addr[1560] = 746;
        test_data[1560] = 33'd2402779610;
        test_addr[1561] = 747;
        test_data[1561] = 33'd4029219969;
        test_addr[1562] = 478;
        test_data[1562] = 33'd6683785524;
        test_addr[1563] = 479;
        test_data[1563] = 33'd271749932;
        test_addr[1564] = 480;
        test_data[1564] = 33'd6399028398;
        test_addr[1565] = 481;
        test_data[1565] = 33'd4465638756;
        test_addr[1566] = 482;
        test_data[1566] = 33'd5003911412;
        test_addr[1567] = 483;
        test_data[1567] = 33'd7895859579;
        test_addr[1568] = 748;
        test_data[1568] = 33'd1620627030;
        test_addr[1569] = 259;
        test_data[1569] = 33'd6361774264;
        test_addr[1570] = 260;
        test_data[1570] = 33'd3784376997;
        test_addr[1571] = 261;
        test_data[1571] = 33'd5923090146;
        test_addr[1572] = 262;
        test_data[1572] = 33'd8172019734;
        test_addr[1573] = 263;
        test_data[1573] = 33'd1168259603;
        test_addr[1574] = 264;
        test_data[1574] = 33'd3017312274;
        test_addr[1575] = 265;
        test_data[1575] = 33'd4232753553;
        test_addr[1576] = 749;
        test_data[1576] = 33'd428043726;
        test_addr[1577] = 750;
        test_data[1577] = 33'd7346017081;
        test_addr[1578] = 234;
        test_data[1578] = 33'd2569948806;
        test_addr[1579] = 235;
        test_data[1579] = 33'd2173127971;
        test_addr[1580] = 236;
        test_data[1580] = 33'd543005921;
        test_addr[1581] = 237;
        test_data[1581] = 33'd2163671273;
        test_addr[1582] = 238;
        test_data[1582] = 33'd1309914105;
        test_addr[1583] = 239;
        test_data[1583] = 33'd6402864615;
        test_addr[1584] = 240;
        test_data[1584] = 33'd1564295992;
        test_addr[1585] = 241;
        test_data[1585] = 33'd5133706534;
        test_addr[1586] = 242;
        test_data[1586] = 33'd6470928813;
        test_addr[1587] = 243;
        test_data[1587] = 33'd3695880751;
        test_addr[1588] = 244;
        test_data[1588] = 33'd3986444448;
        test_addr[1589] = 245;
        test_data[1589] = 33'd2800396312;
        test_addr[1590] = 246;
        test_data[1590] = 33'd2440705799;
        test_addr[1591] = 247;
        test_data[1591] = 33'd8576053712;
        test_addr[1592] = 248;
        test_data[1592] = 33'd2335357878;
        test_addr[1593] = 249;
        test_data[1593] = 33'd1002837958;
        test_addr[1594] = 250;
        test_data[1594] = 33'd2580201917;
        test_addr[1595] = 251;
        test_data[1595] = 33'd1827628710;
        test_addr[1596] = 252;
        test_data[1596] = 33'd2539467430;
        test_addr[1597] = 253;
        test_data[1597] = 33'd1046892784;
        test_addr[1598] = 254;
        test_data[1598] = 33'd893686890;
        test_addr[1599] = 751;
        test_data[1599] = 33'd500787216;
        test_addr[1600] = 148;
        test_data[1600] = 33'd1327006217;
        test_addr[1601] = 149;
        test_data[1601] = 33'd1476414796;
        test_addr[1602] = 150;
        test_data[1602] = 33'd2726814038;
        test_addr[1603] = 151;
        test_data[1603] = 33'd232230619;
        test_addr[1604] = 152;
        test_data[1604] = 33'd7011411635;
        test_addr[1605] = 153;
        test_data[1605] = 33'd5222639249;
        test_addr[1606] = 154;
        test_data[1606] = 33'd6180212131;
        test_addr[1607] = 155;
        test_data[1607] = 33'd1633875019;
        test_addr[1608] = 752;
        test_data[1608] = 33'd5741642759;
        test_addr[1609] = 753;
        test_data[1609] = 33'd3199516579;
        test_addr[1610] = 754;
        test_data[1610] = 33'd733598019;
        test_addr[1611] = 755;
        test_data[1611] = 33'd3037275798;
        test_addr[1612] = 343;
        test_data[1612] = 33'd3938949624;
        test_addr[1613] = 344;
        test_data[1613] = 33'd7588298377;
        test_addr[1614] = 756;
        test_data[1614] = 33'd943611231;
        test_addr[1615] = 757;
        test_data[1615] = 33'd2785722476;
        test_addr[1616] = 758;
        test_data[1616] = 33'd848987015;
        test_addr[1617] = 759;
        test_data[1617] = 33'd8360934625;
        test_addr[1618] = 760;
        test_data[1618] = 33'd5493616857;
        test_addr[1619] = 761;
        test_data[1619] = 33'd1930378489;
        test_addr[1620] = 762;
        test_data[1620] = 33'd8362440394;
        test_addr[1621] = 763;
        test_data[1621] = 33'd3670633852;
        test_addr[1622] = 764;
        test_data[1622] = 33'd5077797580;
        test_addr[1623] = 187;
        test_data[1623] = 33'd6617346832;
        test_addr[1624] = 188;
        test_data[1624] = 33'd3828919794;
        test_addr[1625] = 189;
        test_data[1625] = 33'd2152553771;
        test_addr[1626] = 190;
        test_data[1626] = 33'd7181094638;
        test_addr[1627] = 191;
        test_data[1627] = 33'd1659134554;
        test_addr[1628] = 192;
        test_data[1628] = 33'd323437583;
        test_addr[1629] = 193;
        test_data[1629] = 33'd1908158991;
        test_addr[1630] = 194;
        test_data[1630] = 33'd5817126030;
        test_addr[1631] = 195;
        test_data[1631] = 33'd3019549800;
        test_addr[1632] = 196;
        test_data[1632] = 33'd3889204301;
        test_addr[1633] = 197;
        test_data[1633] = 33'd5108767104;
        test_addr[1634] = 198;
        test_data[1634] = 33'd400801465;
        test_addr[1635] = 199;
        test_data[1635] = 33'd3992018582;
        test_addr[1636] = 200;
        test_data[1636] = 33'd3223549335;
        test_addr[1637] = 201;
        test_data[1637] = 33'd2012336102;
        test_addr[1638] = 202;
        test_data[1638] = 33'd5465287200;
        test_addr[1639] = 203;
        test_data[1639] = 33'd2685333552;
        test_addr[1640] = 204;
        test_data[1640] = 33'd3227643862;
        test_addr[1641] = 205;
        test_data[1641] = 33'd540360476;
        test_addr[1642] = 206;
        test_data[1642] = 33'd2946247101;
        test_addr[1643] = 207;
        test_data[1643] = 33'd5663469898;
        test_addr[1644] = 208;
        test_data[1644] = 33'd1843892378;
        test_addr[1645] = 209;
        test_data[1645] = 33'd5093141273;
        test_addr[1646] = 210;
        test_data[1646] = 33'd6291525726;
        test_addr[1647] = 211;
        test_data[1647] = 33'd3948687695;
        test_addr[1648] = 212;
        test_data[1648] = 33'd3897575557;
        test_addr[1649] = 213;
        test_data[1649] = 33'd1862765609;
        test_addr[1650] = 214;
        test_data[1650] = 33'd3563881117;
        test_addr[1651] = 215;
        test_data[1651] = 33'd584436490;
        test_addr[1652] = 216;
        test_data[1652] = 33'd313568208;
        test_addr[1653] = 217;
        test_data[1653] = 33'd2173355106;
        test_addr[1654] = 218;
        test_data[1654] = 33'd3295815568;
        test_addr[1655] = 219;
        test_data[1655] = 33'd1970268263;
        test_addr[1656] = 220;
        test_data[1656] = 33'd3319839920;
        test_addr[1657] = 221;
        test_data[1657] = 33'd6462431575;
        test_addr[1658] = 222;
        test_data[1658] = 33'd2498690093;
        test_addr[1659] = 223;
        test_data[1659] = 33'd5098110190;
        test_addr[1660] = 224;
        test_data[1660] = 33'd8811210;
        test_addr[1661] = 225;
        test_data[1661] = 33'd6956261276;
        test_addr[1662] = 226;
        test_data[1662] = 33'd2431492093;
        test_addr[1663] = 227;
        test_data[1663] = 33'd4109066461;
        test_addr[1664] = 228;
        test_data[1664] = 33'd4951133192;
        test_addr[1665] = 229;
        test_data[1665] = 33'd2383148880;
        test_addr[1666] = 765;
        test_data[1666] = 33'd6654335476;
        test_addr[1667] = 766;
        test_data[1667] = 33'd1936387940;
        test_addr[1668] = 580;
        test_data[1668] = 33'd4533915551;
        test_addr[1669] = 581;
        test_data[1669] = 33'd7903122207;
        test_addr[1670] = 582;
        test_data[1670] = 33'd3828164037;
        test_addr[1671] = 583;
        test_data[1671] = 33'd5243732807;
        test_addr[1672] = 584;
        test_data[1672] = 33'd3190759241;
        test_addr[1673] = 585;
        test_data[1673] = 33'd6347755539;
        test_addr[1674] = 767;
        test_data[1674] = 33'd1779844196;
        test_addr[1675] = 768;
        test_data[1675] = 33'd3269737958;
        test_addr[1676] = 769;
        test_data[1676] = 33'd7966498928;
        test_addr[1677] = 770;
        test_data[1677] = 33'd2728342669;
        test_addr[1678] = 504;
        test_data[1678] = 33'd2260143172;
        test_addr[1679] = 505;
        test_data[1679] = 33'd4645730717;
        test_addr[1680] = 506;
        test_data[1680] = 33'd4288738455;
        test_addr[1681] = 507;
        test_data[1681] = 33'd6041917015;
        test_addr[1682] = 508;
        test_data[1682] = 33'd1676312471;
        test_addr[1683] = 509;
        test_data[1683] = 33'd4840481955;
        test_addr[1684] = 510;
        test_data[1684] = 33'd6478663792;
        test_addr[1685] = 511;
        test_data[1685] = 33'd1421325492;
        test_addr[1686] = 771;
        test_data[1686] = 33'd2140434203;
        test_addr[1687] = 772;
        test_data[1687] = 33'd2174708313;
        test_addr[1688] = 773;
        test_data[1688] = 33'd5145560188;
        test_addr[1689] = 774;
        test_data[1689] = 33'd773021249;
        test_addr[1690] = 775;
        test_data[1690] = 33'd193689677;
        test_addr[1691] = 776;
        test_data[1691] = 33'd2103915868;
        test_addr[1692] = 777;
        test_data[1692] = 33'd3351668101;
        test_addr[1693] = 778;
        test_data[1693] = 33'd1485151742;
        test_addr[1694] = 779;
        test_data[1694] = 33'd25730636;
        test_addr[1695] = 780;
        test_data[1695] = 33'd3449249766;
        test_addr[1696] = 544;
        test_data[1696] = 33'd118999468;
        test_addr[1697] = 545;
        test_data[1697] = 33'd3588739236;
        test_addr[1698] = 546;
        test_data[1698] = 33'd717909476;
        test_addr[1699] = 547;
        test_data[1699] = 33'd1656097789;
        test_addr[1700] = 548;
        test_data[1700] = 33'd3975122350;
        test_addr[1701] = 549;
        test_data[1701] = 33'd5389056239;
        test_addr[1702] = 550;
        test_data[1702] = 33'd5379842447;
        test_addr[1703] = 551;
        test_data[1703] = 33'd3550124624;
        test_addr[1704] = 552;
        test_data[1704] = 33'd1215198203;
        test_addr[1705] = 553;
        test_data[1705] = 33'd1687299562;
        test_addr[1706] = 554;
        test_data[1706] = 33'd1049579336;
        test_addr[1707] = 555;
        test_data[1707] = 33'd2248499919;
        test_addr[1708] = 556;
        test_data[1708] = 33'd2939472687;
        test_addr[1709] = 557;
        test_data[1709] = 33'd985122537;
        test_addr[1710] = 558;
        test_data[1710] = 33'd5206667930;
        test_addr[1711] = 781;
        test_data[1711] = 33'd2618963896;
        test_addr[1712] = 782;
        test_data[1712] = 33'd1895287559;
        test_addr[1713] = 783;
        test_data[1713] = 33'd6443892364;
        test_addr[1714] = 784;
        test_data[1714] = 33'd2409029183;
        test_addr[1715] = 265;
        test_data[1715] = 33'd4232753553;
        test_addr[1716] = 266;
        test_data[1716] = 33'd6058122676;
        test_addr[1717] = 267;
        test_data[1717] = 33'd2666779884;
        test_addr[1718] = 268;
        test_data[1718] = 33'd878985346;
        test_addr[1719] = 785;
        test_data[1719] = 33'd1730244568;
        test_addr[1720] = 786;
        test_data[1720] = 33'd6764646488;
        test_addr[1721] = 787;
        test_data[1721] = 33'd3191758865;
        test_addr[1722] = 512;
        test_data[1722] = 33'd3788029954;
        test_addr[1723] = 513;
        test_data[1723] = 33'd6326321228;
        test_addr[1724] = 514;
        test_data[1724] = 33'd7681610012;
        test_addr[1725] = 515;
        test_data[1725] = 33'd2354318472;
        test_addr[1726] = 516;
        test_data[1726] = 33'd7443370136;
        test_addr[1727] = 517;
        test_data[1727] = 33'd2393872258;
        test_addr[1728] = 518;
        test_data[1728] = 33'd892001372;
        test_addr[1729] = 519;
        test_data[1729] = 33'd705002716;
        test_addr[1730] = 520;
        test_data[1730] = 33'd2190908579;
        test_addr[1731] = 521;
        test_data[1731] = 33'd1306264201;
        test_addr[1732] = 522;
        test_data[1732] = 33'd511760533;
        test_addr[1733] = 523;
        test_data[1733] = 33'd1659053730;
        test_addr[1734] = 524;
        test_data[1734] = 33'd2535488802;
        test_addr[1735] = 525;
        test_data[1735] = 33'd2367555368;
        test_addr[1736] = 526;
        test_data[1736] = 33'd2518142267;
        test_addr[1737] = 788;
        test_data[1737] = 33'd3817033739;
        test_addr[1738] = 789;
        test_data[1738] = 33'd484067223;
        test_addr[1739] = 790;
        test_data[1739] = 33'd1927359054;
        test_addr[1740] = 791;
        test_data[1740] = 33'd4501345682;
        test_addr[1741] = 792;
        test_data[1741] = 33'd8296217759;
        test_addr[1742] = 793;
        test_data[1742] = 33'd1013045164;
        test_addr[1743] = 794;
        test_data[1743] = 33'd1910908914;
        test_addr[1744] = 795;
        test_data[1744] = 33'd2745117317;
        test_addr[1745] = 796;
        test_data[1745] = 33'd3245915395;
        test_addr[1746] = 797;
        test_data[1746] = 33'd757922546;
        test_addr[1747] = 798;
        test_data[1747] = 33'd7379053212;
        test_addr[1748] = 799;
        test_data[1748] = 33'd2115180072;
        test_addr[1749] = 800;
        test_data[1749] = 33'd4736058885;
        test_addr[1750] = 801;
        test_data[1750] = 33'd2873799072;
        test_addr[1751] = 802;
        test_data[1751] = 33'd1922031926;
        test_addr[1752] = 803;
        test_data[1752] = 33'd3660731959;
        test_addr[1753] = 804;
        test_data[1753] = 33'd8171552530;
        test_addr[1754] = 805;
        test_data[1754] = 33'd341095953;
        test_addr[1755] = 806;
        test_data[1755] = 33'd6098749148;
        test_addr[1756] = 847;
        test_data[1756] = 33'd2773855860;
        test_addr[1757] = 848;
        test_data[1757] = 33'd5098290525;
        test_addr[1758] = 849;
        test_data[1758] = 33'd644666857;
        test_addr[1759] = 850;
        test_data[1759] = 33'd3810045984;
        test_addr[1760] = 851;
        test_data[1760] = 33'd1633202550;
        test_addr[1761] = 852;
        test_data[1761] = 33'd3434666825;
        test_addr[1762] = 853;
        test_data[1762] = 33'd564835311;
        test_addr[1763] = 807;
        test_data[1763] = 33'd619472320;
        test_addr[1764] = 808;
        test_data[1764] = 33'd3811340329;
        test_addr[1765] = 809;
        test_data[1765] = 33'd6641337041;
        test_addr[1766] = 810;
        test_data[1766] = 33'd848075204;
        test_addr[1767] = 811;
        test_data[1767] = 33'd1022680166;
        test_addr[1768] = 812;
        test_data[1768] = 33'd8031115319;
        test_addr[1769] = 813;
        test_data[1769] = 33'd6881328782;
        test_addr[1770] = 814;
        test_data[1770] = 33'd7380718950;
        test_addr[1771] = 815;
        test_data[1771] = 33'd8064737349;
        test_addr[1772] = 816;
        test_data[1772] = 33'd1315395646;
        test_addr[1773] = 817;
        test_data[1773] = 33'd788918906;
        test_addr[1774] = 818;
        test_data[1774] = 33'd3877886931;
        test_addr[1775] = 819;
        test_data[1775] = 33'd5829172731;
        test_addr[1776] = 820;
        test_data[1776] = 33'd1595833567;
        test_addr[1777] = 821;
        test_data[1777] = 33'd3943906068;
        test_addr[1778] = 822;
        test_data[1778] = 33'd2522203454;
        test_addr[1779] = 823;
        test_data[1779] = 33'd8513778702;
        test_addr[1780] = 824;
        test_data[1780] = 33'd5643224463;
        test_addr[1781] = 825;
        test_data[1781] = 33'd2605302930;
        test_addr[1782] = 826;
        test_data[1782] = 33'd4533295374;
        test_addr[1783] = 827;
        test_data[1783] = 33'd5950686121;
        test_addr[1784] = 828;
        test_data[1784] = 33'd5926807822;
        test_addr[1785] = 829;
        test_data[1785] = 33'd1668879510;
        test_addr[1786] = 830;
        test_data[1786] = 33'd3958563769;
        test_addr[1787] = 831;
        test_data[1787] = 33'd1616713383;
        test_addr[1788] = 832;
        test_data[1788] = 33'd2891161115;
        test_addr[1789] = 833;
        test_data[1789] = 33'd8206663985;
        test_addr[1790] = 834;
        test_data[1790] = 33'd3031697508;
        test_addr[1791] = 835;
        test_data[1791] = 33'd1986483545;
        test_addr[1792] = 836;
        test_data[1792] = 33'd4946866410;
        test_addr[1793] = 837;
        test_data[1793] = 33'd8154786606;
        test_addr[1794] = 838;
        test_data[1794] = 33'd7919267230;
        test_addr[1795] = 839;
        test_data[1795] = 33'd2174987116;
        test_addr[1796] = 840;
        test_data[1796] = 33'd2773472885;
        test_addr[1797] = 841;
        test_data[1797] = 33'd846659615;
        test_addr[1798] = 842;
        test_data[1798] = 33'd3536331538;
        test_addr[1799] = 843;
        test_data[1799] = 33'd1817785861;
        test_addr[1800] = 844;
        test_data[1800] = 33'd1556922740;
        test_addr[1801] = 845;
        test_data[1801] = 33'd8485802428;
        test_addr[1802] = 846;
        test_data[1802] = 33'd3605947957;
        test_addr[1803] = 847;
        test_data[1803] = 33'd2773855860;
        test_addr[1804] = 848;
        test_data[1804] = 33'd803323229;
        test_addr[1805] = 849;
        test_data[1805] = 33'd644666857;
        test_addr[1806] = 850;
        test_data[1806] = 33'd4966305263;
        test_addr[1807] = 851;
        test_data[1807] = 33'd1633202550;
        test_addr[1808] = 215;
        test_data[1808] = 33'd584436490;
        test_addr[1809] = 216;
        test_data[1809] = 33'd313568208;
        test_addr[1810] = 217;
        test_data[1810] = 33'd2173355106;
        test_addr[1811] = 218;
        test_data[1811] = 33'd3295815568;
        test_addr[1812] = 219;
        test_data[1812] = 33'd1970268263;
        test_addr[1813] = 220;
        test_data[1813] = 33'd5167346619;
        test_addr[1814] = 221;
        test_data[1814] = 33'd2167464279;
        test_addr[1815] = 222;
        test_data[1815] = 33'd4354234312;
        test_addr[1816] = 223;
        test_data[1816] = 33'd7872783413;
        test_addr[1817] = 224;
        test_data[1817] = 33'd5192288545;
        test_addr[1818] = 225;
        test_data[1818] = 33'd5339806532;
        test_addr[1819] = 226;
        test_data[1819] = 33'd2431492093;
        test_addr[1820] = 227;
        test_data[1820] = 33'd4439384531;
        test_addr[1821] = 228;
        test_data[1821] = 33'd7593156462;
        test_addr[1822] = 229;
        test_data[1822] = 33'd8485589287;
        test_addr[1823] = 230;
        test_data[1823] = 33'd5923214538;
        test_addr[1824] = 231;
        test_data[1824] = 33'd1756904191;
        test_addr[1825] = 852;
        test_data[1825] = 33'd3434666825;
        test_addr[1826] = 853;
        test_data[1826] = 33'd564835311;
        test_addr[1827] = 854;
        test_data[1827] = 33'd7225638048;
        test_addr[1828] = 855;
        test_data[1828] = 33'd3981959618;
        test_addr[1829] = 856;
        test_data[1829] = 33'd821321256;
        test_addr[1830] = 857;
        test_data[1830] = 33'd54187291;
        test_addr[1831] = 609;
        test_data[1831] = 33'd7002969478;
        test_addr[1832] = 610;
        test_data[1832] = 33'd2655954426;
        test_addr[1833] = 611;
        test_data[1833] = 33'd507597236;
        test_addr[1834] = 858;
        test_data[1834] = 33'd1198553052;
        test_addr[1835] = 859;
        test_data[1835] = 33'd3073653273;
        test_addr[1836] = 860;
        test_data[1836] = 33'd3552320581;
        test_addr[1837] = 861;
        test_data[1837] = 33'd469402357;
        test_addr[1838] = 862;
        test_data[1838] = 33'd3411959600;
        test_addr[1839] = 863;
        test_data[1839] = 33'd4389617786;
        test_addr[1840] = 864;
        test_data[1840] = 33'd8144291570;
        test_addr[1841] = 95;
        test_data[1841] = 33'd610452162;
        test_addr[1842] = 96;
        test_data[1842] = 33'd3730512133;
        test_addr[1843] = 97;
        test_data[1843] = 33'd654962339;
        test_addr[1844] = 98;
        test_data[1844] = 33'd2789486256;
        test_addr[1845] = 99;
        test_data[1845] = 33'd1718939551;
        test_addr[1846] = 865;
        test_data[1846] = 33'd6443359624;
        test_addr[1847] = 866;
        test_data[1847] = 33'd366355984;
        test_addr[1848] = 701;
        test_data[1848] = 33'd835744670;
        test_addr[1849] = 702;
        test_data[1849] = 33'd1564728561;
        test_addr[1850] = 703;
        test_data[1850] = 33'd1255659046;
        test_addr[1851] = 704;
        test_data[1851] = 33'd5506544236;
        test_addr[1852] = 705;
        test_data[1852] = 33'd1911257944;
        test_addr[1853] = 706;
        test_data[1853] = 33'd3521378079;
        test_addr[1854] = 707;
        test_data[1854] = 33'd3041654547;
        test_addr[1855] = 708;
        test_data[1855] = 33'd3884518045;
        test_addr[1856] = 709;
        test_data[1856] = 33'd3130440955;
        test_addr[1857] = 867;
        test_data[1857] = 33'd8521988990;
        test_addr[1858] = 868;
        test_data[1858] = 33'd5647700588;
        test_addr[1859] = 869;
        test_data[1859] = 33'd5545636895;
        test_addr[1860] = 841;
        test_data[1860] = 33'd6275153422;
        test_addr[1861] = 842;
        test_data[1861] = 33'd3536331538;
        test_addr[1862] = 843;
        test_data[1862] = 33'd1817785861;
        test_addr[1863] = 844;
        test_data[1863] = 33'd7233953608;
        test_addr[1864] = 845;
        test_data[1864] = 33'd4190835132;
        test_addr[1865] = 846;
        test_data[1865] = 33'd3605947957;
        test_addr[1866] = 870;
        test_data[1866] = 33'd8554397087;
        test_addr[1867] = 233;
        test_data[1867] = 33'd1437501823;
        test_addr[1868] = 871;
        test_data[1868] = 33'd4958145258;
        test_addr[1869] = 872;
        test_data[1869] = 33'd7568312576;
        test_addr[1870] = 873;
        test_data[1870] = 33'd2989369719;
        test_addr[1871] = 874;
        test_data[1871] = 33'd7147717618;
        test_addr[1872] = 875;
        test_data[1872] = 33'd4963088180;
        test_addr[1873] = 876;
        test_data[1873] = 33'd4748482911;
        test_addr[1874] = 877;
        test_data[1874] = 33'd1774453158;
        test_addr[1875] = 878;
        test_data[1875] = 33'd1205002421;
        test_addr[1876] = 879;
        test_data[1876] = 33'd2912634867;
        test_addr[1877] = 426;
        test_data[1877] = 33'd3544872180;
        test_addr[1878] = 427;
        test_data[1878] = 33'd6560606145;
        test_addr[1879] = 428;
        test_data[1879] = 33'd4592660939;
        test_addr[1880] = 429;
        test_data[1880] = 33'd4250490692;
        test_addr[1881] = 430;
        test_data[1881] = 33'd4300700850;
        test_addr[1882] = 431;
        test_data[1882] = 33'd2790016042;
        test_addr[1883] = 432;
        test_data[1883] = 33'd3691339593;
        test_addr[1884] = 433;
        test_data[1884] = 33'd1999264964;
        test_addr[1885] = 434;
        test_data[1885] = 33'd5959374967;
        test_addr[1886] = 880;
        test_data[1886] = 33'd2614693622;
        test_addr[1887] = 881;
        test_data[1887] = 33'd4981615445;
        test_addr[1888] = 882;
        test_data[1888] = 33'd809342124;
        test_addr[1889] = 883;
        test_data[1889] = 33'd997878904;
        test_addr[1890] = 884;
        test_data[1890] = 33'd665306548;
        test_addr[1891] = 885;
        test_data[1891] = 33'd6252126588;
        test_addr[1892] = 886;
        test_data[1892] = 33'd7893206211;
        test_addr[1893] = 887;
        test_data[1893] = 33'd2450826475;
        test_addr[1894] = 394;
        test_data[1894] = 33'd7935146232;
        test_addr[1895] = 888;
        test_data[1895] = 33'd7610999202;
        test_addr[1896] = 889;
        test_data[1896] = 33'd858761786;
        test_addr[1897] = 890;
        test_data[1897] = 33'd3932332099;
        test_addr[1898] = 891;
        test_data[1898] = 33'd1541522239;
        test_addr[1899] = 676;
        test_data[1899] = 33'd1104785019;
        test_addr[1900] = 677;
        test_data[1900] = 33'd929867826;
        test_addr[1901] = 678;
        test_data[1901] = 33'd1236351052;
        test_addr[1902] = 679;
        test_data[1902] = 33'd8102253042;
        test_addr[1903] = 680;
        test_data[1903] = 33'd3119041072;
        test_addr[1904] = 892;
        test_data[1904] = 33'd7635632030;
        test_addr[1905] = 893;
        test_data[1905] = 33'd7392298970;
        test_addr[1906] = 894;
        test_data[1906] = 33'd1045852187;
        test_addr[1907] = 895;
        test_data[1907] = 33'd119509833;
        test_addr[1908] = 896;
        test_data[1908] = 33'd298321624;
        test_addr[1909] = 941;
        test_data[1909] = 33'd2633217852;
        test_addr[1910] = 942;
        test_data[1910] = 33'd2811349348;
        test_addr[1911] = 897;
        test_data[1911] = 33'd2281912767;
        test_addr[1912] = 898;
        test_data[1912] = 33'd262579741;
        test_addr[1913] = 899;
        test_data[1913] = 33'd3207744075;
        test_addr[1914] = 900;
        test_data[1914] = 33'd3651982289;
        test_addr[1915] = 901;
        test_data[1915] = 33'd1575034248;
        test_addr[1916] = 902;
        test_data[1916] = 33'd910704321;
        test_addr[1917] = 903;
        test_data[1917] = 33'd4562001145;
        test_addr[1918] = 904;
        test_data[1918] = 33'd2673042208;
        test_addr[1919] = 905;
        test_data[1919] = 33'd8329224496;
        test_addr[1920] = 906;
        test_data[1920] = 33'd774256557;
        test_addr[1921] = 907;
        test_data[1921] = 33'd901261549;
        test_addr[1922] = 908;
        test_data[1922] = 33'd2319053902;
        test_addr[1923] = 909;
        test_data[1923] = 33'd1962590118;
        test_addr[1924] = 910;
        test_data[1924] = 33'd885454967;
        test_addr[1925] = 911;
        test_data[1925] = 33'd5274849057;
        test_addr[1926] = 912;
        test_data[1926] = 33'd7536609840;
        test_addr[1927] = 913;
        test_data[1927] = 33'd3108154670;
        test_addr[1928] = 914;
        test_data[1928] = 33'd4329753202;
        test_addr[1929] = 915;
        test_data[1929] = 33'd1563133648;
        test_addr[1930] = 916;
        test_data[1930] = 33'd4396484440;
        test_addr[1931] = 917;
        test_data[1931] = 33'd4071938350;
        test_addr[1932] = 918;
        test_data[1932] = 33'd5073500082;
        test_addr[1933] = 919;
        test_data[1933] = 33'd7402224095;
        test_addr[1934] = 920;
        test_data[1934] = 33'd3915123610;
        test_addr[1935] = 921;
        test_data[1935] = 33'd5539980728;
        test_addr[1936] = 922;
        test_data[1936] = 33'd5414210260;
        test_addr[1937] = 879;
        test_data[1937] = 33'd4961280741;
        test_addr[1938] = 880;
        test_data[1938] = 33'd2614693622;
        test_addr[1939] = 881;
        test_data[1939] = 33'd686648149;
        test_addr[1940] = 882;
        test_data[1940] = 33'd8256080387;
        test_addr[1941] = 923;
        test_data[1941] = 33'd7398512428;
        test_addr[1942] = 924;
        test_data[1942] = 33'd5888758377;
        test_addr[1943] = 925;
        test_data[1943] = 33'd1313195782;
        test_addr[1944] = 926;
        test_data[1944] = 33'd4642543402;
        test_addr[1945] = 927;
        test_data[1945] = 33'd8562606539;
        test_addr[1946] = 928;
        test_data[1946] = 33'd5389355337;
        test_addr[1947] = 929;
        test_data[1947] = 33'd1467497009;
        test_addr[1948] = 930;
        test_data[1948] = 33'd1729249679;
        test_addr[1949] = 931;
        test_data[1949] = 33'd1776715744;
        test_addr[1950] = 932;
        test_data[1950] = 33'd360085129;
        test_addr[1951] = 933;
        test_data[1951] = 33'd4810103766;
        test_addr[1952] = 934;
        test_data[1952] = 33'd392045396;
        test_addr[1953] = 935;
        test_data[1953] = 33'd2632191667;
        test_addr[1954] = 936;
        test_data[1954] = 33'd3408512394;
        test_addr[1955] = 937;
        test_data[1955] = 33'd3663858100;
        test_addr[1956] = 938;
        test_data[1956] = 33'd4703518237;
        test_addr[1957] = 939;
        test_data[1957] = 33'd4240778167;
        test_addr[1958] = 940;
        test_data[1958] = 33'd338549878;
        test_addr[1959] = 941;
        test_data[1959] = 33'd7506804988;
        test_addr[1960] = 942;
        test_data[1960] = 33'd5214716528;
        test_addr[1961] = 943;
        test_data[1961] = 33'd5305954539;
        test_addr[1962] = 944;
        test_data[1962] = 33'd1901157862;
        test_addr[1963] = 945;
        test_data[1963] = 33'd4453432581;
        test_addr[1964] = 946;
        test_data[1964] = 33'd4251511846;
        test_addr[1965] = 408;
        test_data[1965] = 33'd3784952382;
        test_addr[1966] = 409;
        test_data[1966] = 33'd829691805;
        test_addr[1967] = 410;
        test_data[1967] = 33'd5363043309;
        test_addr[1968] = 411;
        test_data[1968] = 33'd6978074757;
        test_addr[1969] = 412;
        test_data[1969] = 33'd1038301027;
        test_addr[1970] = 413;
        test_data[1970] = 33'd2856665508;
        test_addr[1971] = 414;
        test_data[1971] = 33'd8539748194;
        test_addr[1972] = 415;
        test_data[1972] = 33'd268942874;
        test_addr[1973] = 416;
        test_data[1973] = 33'd2315947450;
        test_addr[1974] = 417;
        test_data[1974] = 33'd2168180925;
        test_addr[1975] = 418;
        test_data[1975] = 33'd3119127120;
        test_addr[1976] = 419;
        test_data[1976] = 33'd3511401386;
        test_addr[1977] = 420;
        test_data[1977] = 33'd6963080496;
        test_addr[1978] = 421;
        test_data[1978] = 33'd257964552;
        test_addr[1979] = 422;
        test_data[1979] = 33'd962672775;
        test_addr[1980] = 423;
        test_data[1980] = 33'd3728980285;
        test_addr[1981] = 424;
        test_data[1981] = 33'd5485871675;
        test_addr[1982] = 425;
        test_data[1982] = 33'd3494559305;
        test_addr[1983] = 426;
        test_data[1983] = 33'd3544872180;
        test_addr[1984] = 427;
        test_data[1984] = 33'd2265638849;
        test_addr[1985] = 428;
        test_data[1985] = 33'd4686255400;
        test_addr[1986] = 429;
        test_data[1986] = 33'd6477767881;
        test_addr[1987] = 947;
        test_data[1987] = 33'd6085266752;
        test_addr[1988] = 948;
        test_data[1988] = 33'd4990492510;
        test_addr[1989] = 949;
        test_data[1989] = 33'd525044368;
        test_addr[1990] = 950;
        test_data[1990] = 33'd2680314078;
        test_addr[1991] = 951;
        test_data[1991] = 33'd2339532244;
        test_addr[1992] = 952;
        test_data[1992] = 33'd4040559479;
        test_addr[1993] = 953;
        test_data[1993] = 33'd8187851353;
        test_addr[1994] = 954;
        test_data[1994] = 33'd920008339;
        test_addr[1995] = 955;
        test_data[1995] = 33'd6454584696;
        test_addr[1996] = 956;
        test_data[1996] = 33'd922515263;
        test_addr[1997] = 893;
        test_data[1997] = 33'd3097331674;
        test_addr[1998] = 894;
        test_data[1998] = 33'd1045852187;
        test_addr[1999] = 895;
        test_data[1999] = 33'd5770680254;
        test_addr[2000] = 896;
        test_data[2000] = 33'd8369082223;
        test_addr[2001] = 897;
        test_data[2001] = 33'd4966421913;
        test_addr[2002] = 898;
        test_data[2002] = 33'd262579741;
        test_addr[2003] = 899;
        test_data[2003] = 33'd3207744075;
        test_addr[2004] = 900;
        test_data[2004] = 33'd4892274530;
        test_addr[2005] = 901;
        test_data[2005] = 33'd6137988933;
        test_addr[2006] = 902;
        test_data[2006] = 33'd910704321;
        test_addr[2007] = 903;
        test_data[2007] = 33'd267033849;
        test_addr[2008] = 904;
        test_data[2008] = 33'd2673042208;
        test_addr[2009] = 905;
        test_data[2009] = 33'd4034257200;
        test_addr[2010] = 906;
        test_data[2010] = 33'd774256557;
        test_addr[2011] = 907;
        test_data[2011] = 33'd901261549;
        test_addr[2012] = 908;
        test_data[2012] = 33'd2319053902;
        test_addr[2013] = 909;
        test_data[2013] = 33'd1962590118;
        test_addr[2014] = 910;
        test_data[2014] = 33'd7194778027;
        test_addr[2015] = 911;
        test_data[2015] = 33'd7400768278;
        test_addr[2016] = 912;
        test_data[2016] = 33'd3241642544;
        test_addr[2017] = 913;
        test_data[2017] = 33'd6536880563;
        test_addr[2018] = 957;
        test_data[2018] = 33'd8020902385;
        test_addr[2019] = 174;
        test_data[2019] = 33'd4464925744;
        test_addr[2020] = 175;
        test_data[2020] = 33'd1951074742;
        test_addr[2021] = 176;
        test_data[2021] = 33'd6718116146;
        test_addr[2022] = 177;
        test_data[2022] = 33'd2547298871;
        test_addr[2023] = 178;
        test_data[2023] = 33'd1390194371;
        test_addr[2024] = 958;
        test_data[2024] = 33'd1131678623;
        test_addr[2025] = 959;
        test_data[2025] = 33'd3011059689;
        test_addr[2026] = 960;
        test_data[2026] = 33'd813414639;
        test_addr[2027] = 961;
        test_data[2027] = 33'd2648618923;
        test_addr[2028] = 970;
        test_data[2028] = 33'd1523162636;
        test_addr[2029] = 971;
        test_data[2029] = 33'd1160760996;
        test_addr[2030] = 972;
        test_data[2030] = 33'd764522856;
        test_addr[2031] = 973;
        test_data[2031] = 33'd5401070589;
        test_addr[2032] = 974;
        test_data[2032] = 33'd5145408456;
        test_addr[2033] = 975;
        test_data[2033] = 33'd902628290;
        test_addr[2034] = 976;
        test_data[2034] = 33'd7814211820;
        test_addr[2035] = 977;
        test_data[2035] = 33'd275231142;
        test_addr[2036] = 962;
        test_data[2036] = 33'd3660914740;
        test_addr[2037] = 963;
        test_data[2037] = 33'd3778906056;
        test_addr[2038] = 964;
        test_data[2038] = 33'd1676243570;
        test_addr[2039] = 965;
        test_data[2039] = 33'd533232901;
        test_addr[2040] = 794;
        test_data[2040] = 33'd1910908914;
        test_addr[2041] = 795;
        test_data[2041] = 33'd2745117317;
        test_addr[2042] = 796;
        test_data[2042] = 33'd3245915395;
        test_addr[2043] = 797;
        test_data[2043] = 33'd757922546;
        test_addr[2044] = 798;
        test_data[2044] = 33'd3084085916;
        test_addr[2045] = 799;
        test_data[2045] = 33'd2115180072;
        test_addr[2046] = 800;
        test_data[2046] = 33'd6750953126;
        test_addr[2047] = 801;
        test_data[2047] = 33'd2873799072;
        test_addr[2048] = 802;
        test_data[2048] = 33'd1922031926;
        test_addr[2049] = 803;
        test_data[2049] = 33'd3660731959;
        test_addr[2050] = 804;
        test_data[2050] = 33'd3876585234;
        test_addr[2051] = 805;
        test_data[2051] = 33'd341095953;
        test_addr[2052] = 966;
        test_data[2052] = 33'd4814917696;
        test_addr[2053] = 967;
        test_data[2053] = 33'd2540554632;
        test_addr[2054] = 297;
        test_data[2054] = 33'd3121280700;
        test_addr[2055] = 298;
        test_data[2055] = 33'd7287873986;
        test_addr[2056] = 299;
        test_data[2056] = 33'd7925509197;
        test_addr[2057] = 300;
        test_data[2057] = 33'd1786211448;
        test_addr[2058] = 301;
        test_data[2058] = 33'd178124090;
        test_addr[2059] = 302;
        test_data[2059] = 33'd3250392161;
        test_addr[2060] = 303;
        test_data[2060] = 33'd4613104053;
        test_addr[2061] = 304;
        test_data[2061] = 33'd8222582424;
        test_addr[2062] = 305;
        test_data[2062] = 33'd6291057851;
        test_addr[2063] = 306;
        test_data[2063] = 33'd8366320762;
        test_addr[2064] = 968;
        test_data[2064] = 33'd759450314;
        test_addr[2065] = 969;
        test_data[2065] = 33'd4246657183;
        test_addr[2066] = 970;
        test_data[2066] = 33'd1523162636;
        test_addr[2067] = 971;
        test_data[2067] = 33'd1160760996;
        test_addr[2068] = 972;
        test_data[2068] = 33'd764522856;
        test_addr[2069] = 973;
        test_data[2069] = 33'd1106103293;
        test_addr[2070] = 974;
        test_data[2070] = 33'd8132737090;
        test_addr[2071] = 975;
        test_data[2071] = 33'd8178522233;
        test_addr[2072] = 976;
        test_data[2072] = 33'd3519244524;
        test_addr[2073] = 977;
        test_data[2073] = 33'd275231142;
        test_addr[2074] = 978;
        test_data[2074] = 33'd2338947152;
        test_addr[2075] = 979;
        test_data[2075] = 33'd4378473381;
        test_addr[2076] = 980;
        test_data[2076] = 33'd2034359482;
        test_addr[2077] = 981;
        test_data[2077] = 33'd318233107;
        test_addr[2078] = 982;
        test_data[2078] = 33'd4040828699;
        test_addr[2079] = 983;
        test_data[2079] = 33'd1211923792;
        test_addr[2080] = 71;
        test_data[2080] = 33'd7369205226;
        test_addr[2081] = 72;
        test_data[2081] = 33'd7031374970;
        test_addr[2082] = 73;
        test_data[2082] = 33'd1855683855;
        test_addr[2083] = 984;
        test_data[2083] = 33'd2842558085;
        test_addr[2084] = 985;
        test_data[2084] = 33'd6141540249;
        test_addr[2085] = 986;
        test_data[2085] = 33'd4830666324;
        test_addr[2086] = 987;
        test_data[2086] = 33'd3038027771;
        test_addr[2087] = 988;
        test_data[2087] = 33'd271887483;
        test_addr[2088] = 989;
        test_data[2088] = 33'd2221065516;
        test_addr[2089] = 441;
        test_data[2089] = 33'd7847970210;
        test_addr[2090] = 442;
        test_data[2090] = 33'd2891047966;
        test_addr[2091] = 443;
        test_data[2091] = 33'd7027893677;
        test_addr[2092] = 990;
        test_data[2092] = 33'd3379643487;
        test_addr[2093] = 991;
        test_data[2093] = 33'd2418675797;
        test_addr[2094] = 992;
        test_data[2094] = 33'd964179193;
        test_addr[2095] = 210;
        test_data[2095] = 33'd1996558430;
        test_addr[2096] = 211;
        test_data[2096] = 33'd3948687695;
        test_addr[2097] = 993;
        test_data[2097] = 33'd8493614423;
        test_addr[2098] = 994;
        test_data[2098] = 33'd2733544077;
        test_addr[2099] = 995;
        test_data[2099] = 33'd3745988993;
        test_addr[2100] = 996;
        test_data[2100] = 33'd6923613209;
        test_addr[2101] = 997;
        test_data[2101] = 33'd1759334156;
        test_addr[2102] = 998;
        test_data[2102] = 33'd1827708917;
        test_addr[2103] = 999;
        test_data[2103] = 33'd2104347660;
        test_addr[2104] = 1000;
        test_data[2104] = 33'd116060540;
        test_addr[2105] = 1001;
        test_data[2105] = 33'd4495122067;
        test_addr[2106] = 1002;
        test_data[2106] = 33'd8209930010;
        test_addr[2107] = 870;
        test_data[2107] = 33'd4259429791;
        test_addr[2108] = 871;
        test_data[2108] = 33'd8414268803;
        test_addr[2109] = 872;
        test_data[2109] = 33'd4857656037;
        test_addr[2110] = 873;
        test_data[2110] = 33'd4480685481;
        test_addr[2111] = 874;
        test_data[2111] = 33'd2852750322;
        test_addr[2112] = 875;
        test_data[2112] = 33'd668120884;
        test_addr[2113] = 1003;
        test_data[2113] = 33'd5085340007;
        test_addr[2114] = 1004;
        test_data[2114] = 33'd2099492465;
        test_addr[2115] = 1005;
        test_data[2115] = 33'd4830371818;
        test_addr[2116] = 1006;
        test_data[2116] = 33'd7683870550;
        test_addr[2117] = 1007;
        test_data[2117] = 33'd166563627;
        test_addr[2118] = 1008;
        test_data[2118] = 33'd4215858546;
        test_addr[2119] = 1009;
        test_data[2119] = 33'd1316389492;
        test_addr[2120] = 938;
        test_data[2120] = 33'd408550941;
        test_addr[2121] = 939;
        test_data[2121] = 33'd5462751640;
        test_addr[2122] = 940;
        test_data[2122] = 33'd7522727880;
        test_addr[2123] = 941;
        test_data[2123] = 33'd8486645090;
        test_addr[2124] = 942;
        test_data[2124] = 33'd919749232;
        test_addr[2125] = 943;
        test_data[2125] = 33'd1010987243;
        test_addr[2126] = 1010;
        test_data[2126] = 33'd3511528593;
        test_addr[2127] = 160;
        test_data[2127] = 33'd2802001540;
        test_addr[2128] = 161;
        test_data[2128] = 33'd260760954;
        test_addr[2129] = 162;
        test_data[2129] = 33'd760186910;
        test_addr[2130] = 163;
        test_data[2130] = 33'd5506713493;
        test_addr[2131] = 164;
        test_data[2131] = 33'd3847429411;
        test_addr[2132] = 1011;
        test_data[2132] = 33'd133678878;
        test_addr[2133] = 172;
        test_data[2133] = 33'd5351356825;
        test_addr[2134] = 173;
        test_data[2134] = 33'd6197345921;
        test_addr[2135] = 174;
        test_data[2135] = 33'd169958448;
        test_addr[2136] = 175;
        test_data[2136] = 33'd1951074742;
        test_addr[2137] = 176;
        test_data[2137] = 33'd7132708773;
        test_addr[2138] = 177;
        test_data[2138] = 33'd2547298871;
        test_addr[2139] = 178;
        test_data[2139] = 33'd1390194371;
        test_addr[2140] = 1012;
        test_data[2140] = 33'd1486798971;
        test_addr[2141] = 1013;
        test_data[2141] = 33'd7338791364;
        test_addr[2142] = 1014;
        test_data[2142] = 33'd5434081504;
        test_addr[2143] = 1015;
        test_data[2143] = 33'd4466770648;
        test_addr[2144] = 1016;
        test_data[2144] = 33'd2042201759;
        test_addr[2145] = 1017;
        test_data[2145] = 33'd4871860239;
        test_addr[2146] = 1018;
        test_data[2146] = 33'd2984861369;
        test_addr[2147] = 1019;
        test_data[2147] = 33'd5665402705;
        test_addr[2148] = 1020;
        test_data[2148] = 33'd5956439698;
        test_addr[2149] = 1021;
        test_data[2149] = 33'd229156893;
        test_addr[2150] = 1022;
        test_data[2150] = 33'd657762763;
        test_addr[2151] = 586;
        test_data[2151] = 33'd3389351130;
        test_addr[2152] = 587;
        test_data[2152] = 33'd4511711526;
        test_addr[2153] = 588;
        test_data[2153] = 33'd7871883137;
        test_addr[2154] = 589;
        test_data[2154] = 33'd7614033787;
        test_addr[2155] = 590;
        test_data[2155] = 33'd8412362183;
        test_addr[2156] = 591;
        test_data[2156] = 33'd3818804376;
        test_addr[2157] = 592;
        test_data[2157] = 33'd5275653564;
        test_addr[2158] = 593;
        test_data[2158] = 33'd4098723952;
        test_addr[2159] = 594;
        test_data[2159] = 33'd2232370504;
        test_addr[2160] = 595;
        test_data[2160] = 33'd7968629194;
        test_addr[2161] = 596;
        test_data[2161] = 33'd3894227902;
        test_addr[2162] = 597;
        test_data[2162] = 33'd6684693016;
        test_addr[2163] = 598;
        test_data[2163] = 33'd133191090;
        test_addr[2164] = 599;
        test_data[2164] = 33'd2221731456;
        test_addr[2165] = 600;
        test_data[2165] = 33'd2084621993;
        test_addr[2166] = 601;
        test_data[2166] = 33'd1528966083;
        test_addr[2167] = 602;
        test_data[2167] = 33'd2985258556;
        test_addr[2168] = 603;
        test_data[2168] = 33'd1521945037;
        test_addr[2169] = 604;
        test_data[2169] = 33'd2543781384;
        test_addr[2170] = 605;
        test_data[2170] = 33'd2631117550;
        test_addr[2171] = 606;
        test_data[2171] = 33'd318066958;
        test_addr[2172] = 1023;
        test_data[2172] = 33'd2095860060;
        test_addr[2173] = 0;
        test_data[2173] = 33'd597582581;
        test_addr[2174] = 1;
        test_data[2174] = 33'd4660195457;
        test_addr[2175] = 2;
        test_data[2175] = 33'd244488320;
        test_addr[2176] = 3;
        test_data[2176] = 33'd2009627834;
        test_addr[2177] = 4;
        test_data[2177] = 33'd1187404859;
        test_addr[2178] = 5;
        test_data[2178] = 33'd6841050661;
        test_addr[2179] = 6;
        test_data[2179] = 33'd3021698007;
        test_addr[2180] = 7;
        test_data[2180] = 33'd8317924608;
        test_addr[2181] = 8;
        test_data[2181] = 33'd4074274575;
        test_addr[2182] = 831;
        test_data[2182] = 33'd4459705183;
        test_addr[2183] = 832;
        test_data[2183] = 33'd2891161115;
        test_addr[2184] = 833;
        test_data[2184] = 33'd3911696689;
        test_addr[2185] = 834;
        test_data[2185] = 33'd7705026509;
        test_addr[2186] = 835;
        test_data[2186] = 33'd7359431071;
        test_addr[2187] = 836;
        test_data[2187] = 33'd651899114;
        test_addr[2188] = 9;
        test_data[2188] = 33'd2158628397;
        test_addr[2189] = 10;
        test_data[2189] = 33'd2770097472;
        test_addr[2190] = 444;
        test_data[2190] = 33'd2972090766;
        test_addr[2191] = 445;
        test_data[2191] = 33'd2392101323;
        test_addr[2192] = 446;
        test_data[2192] = 33'd7276178833;
        test_addr[2193] = 447;
        test_data[2193] = 33'd1470049012;
        test_addr[2194] = 448;
        test_data[2194] = 33'd4639034570;
        test_addr[2195] = 449;
        test_data[2195] = 33'd557852968;
        test_addr[2196] = 450;
        test_data[2196] = 33'd5826480136;
        test_addr[2197] = 451;
        test_data[2197] = 33'd1824370581;
        test_addr[2198] = 452;
        test_data[2198] = 33'd1349213303;
        test_addr[2199] = 453;
        test_data[2199] = 33'd4417027083;
        test_addr[2200] = 454;
        test_data[2200] = 33'd3918291114;
        test_addr[2201] = 455;
        test_data[2201] = 33'd1395496028;
        test_addr[2202] = 456;
        test_data[2202] = 33'd3486845368;
        test_addr[2203] = 457;
        test_data[2203] = 33'd5639993044;
        test_addr[2204] = 458;
        test_data[2204] = 33'd833450510;
        test_addr[2205] = 459;
        test_data[2205] = 33'd826235681;
        test_addr[2206] = 460;
        test_data[2206] = 33'd3390313948;
        test_addr[2207] = 461;
        test_data[2207] = 33'd1580710012;
        test_addr[2208] = 462;
        test_data[2208] = 33'd3770112161;
        test_addr[2209] = 463;
        test_data[2209] = 33'd4010236394;
        test_addr[2210] = 464;
        test_data[2210] = 33'd3147145687;
        test_addr[2211] = 465;
        test_data[2211] = 33'd1076516124;
        test_addr[2212] = 466;
        test_data[2212] = 33'd4780398749;
        test_addr[2213] = 467;
        test_data[2213] = 33'd1263605750;
        test_addr[2214] = 11;
        test_data[2214] = 33'd4191856559;
        test_addr[2215] = 12;
        test_data[2215] = 33'd290304978;
        test_addr[2216] = 13;
        test_data[2216] = 33'd3587268486;
        test_addr[2217] = 14;
        test_data[2217] = 33'd1178385445;
        test_addr[2218] = 15;
        test_data[2218] = 33'd8109089243;
        test_addr[2219] = 16;
        test_data[2219] = 33'd1125683639;
        test_addr[2220] = 17;
        test_data[2220] = 33'd7370988526;
        test_addr[2221] = 18;
        test_data[2221] = 33'd4089621706;
        test_addr[2222] = 19;
        test_data[2222] = 33'd7053565693;
        test_addr[2223] = 20;
        test_data[2223] = 33'd5760168055;
        test_addr[2224] = 21;
        test_data[2224] = 33'd1866610343;
        test_addr[2225] = 876;
        test_data[2225] = 33'd6407374840;
        test_addr[2226] = 877;
        test_data[2226] = 33'd4673563836;
        test_addr[2227] = 878;
        test_data[2227] = 33'd7640490510;
        test_addr[2228] = 879;
        test_data[2228] = 33'd5135258231;
        test_addr[2229] = 880;
        test_data[2229] = 33'd5553403422;
        test_addr[2230] = 22;
        test_data[2230] = 33'd1238017576;
        test_addr[2231] = 23;
        test_data[2231] = 33'd2770618699;
        test_addr[2232] = 24;
        test_data[2232] = 33'd619906137;
        test_addr[2233] = 25;
        test_data[2233] = 33'd3881438871;
        test_addr[2234] = 26;
        test_data[2234] = 33'd7172686920;
        test_addr[2235] = 27;
        test_data[2235] = 33'd2950000704;
        test_addr[2236] = 28;
        test_data[2236] = 33'd2040897048;
        test_addr[2237] = 29;
        test_data[2237] = 33'd580774497;
        test_addr[2238] = 30;
        test_data[2238] = 33'd3252174221;
        test_addr[2239] = 31;
        test_data[2239] = 33'd1738403846;
        test_addr[2240] = 227;
        test_data[2240] = 33'd144417235;
        test_addr[2241] = 228;
        test_data[2241] = 33'd3298189166;
        test_addr[2242] = 229;
        test_data[2242] = 33'd4190621991;
        test_addr[2243] = 230;
        test_data[2243] = 33'd1628247242;
        test_addr[2244] = 231;
        test_data[2244] = 33'd1756904191;
        test_addr[2245] = 232;
        test_data[2245] = 33'd3657253458;
        test_addr[2246] = 233;
        test_data[2246] = 33'd1437501823;
        test_addr[2247] = 234;
        test_data[2247] = 33'd2569948806;
        test_addr[2248] = 235;
        test_data[2248] = 33'd8245569563;
        test_addr[2249] = 236;
        test_data[2249] = 33'd4914842070;
        test_addr[2250] = 237;
        test_data[2250] = 33'd6518665588;
        test_addr[2251] = 238;
        test_data[2251] = 33'd1309914105;
        test_addr[2252] = 239;
        test_data[2252] = 33'd6329125648;
        test_addr[2253] = 240;
        test_data[2253] = 33'd1564295992;
        test_addr[2254] = 241;
        test_data[2254] = 33'd6929919309;
        test_addr[2255] = 242;
        test_data[2255] = 33'd2175961517;
        test_addr[2256] = 243;
        test_data[2256] = 33'd3695880751;
        test_addr[2257] = 244;
        test_data[2257] = 33'd3986444448;
        test_addr[2258] = 245;
        test_data[2258] = 33'd5010090536;
        test_addr[2259] = 246;
        test_data[2259] = 33'd5850686797;
        test_addr[2260] = 32;
        test_data[2260] = 33'd838905011;
        test_addr[2261] = 33;
        test_data[2261] = 33'd1455572206;
        test_addr[2262] = 188;
        test_data[2262] = 33'd7264137225;
        test_addr[2263] = 34;
        test_data[2263] = 33'd3084178052;
        test_addr[2264] = 35;
        test_data[2264] = 33'd273674846;
        test_addr[2265] = 36;
        test_data[2265] = 33'd3086044954;
        test_addr[2266] = 37;
        test_data[2266] = 33'd2005231466;
        test_addr[2267] = 38;
        test_data[2267] = 33'd4009161584;
        test_addr[2268] = 39;
        test_data[2268] = 33'd8566865742;
        test_addr[2269] = 40;
        test_data[2269] = 33'd667246577;
        test_addr[2270] = 41;
        test_data[2270] = 33'd858247705;
        test_addr[2271] = 42;
        test_data[2271] = 33'd7777753368;
        test_addr[2272] = 43;
        test_data[2272] = 33'd8562567809;
        test_addr[2273] = 44;
        test_data[2273] = 33'd7537111177;
        test_addr[2274] = 45;
        test_data[2274] = 33'd1124776585;
        test_addr[2275] = 46;
        test_data[2275] = 33'd6236005639;
        test_addr[2276] = 47;
        test_data[2276] = 33'd167184051;
        test_addr[2277] = 48;
        test_data[2277] = 33'd5447514403;
        test_addr[2278] = 49;
        test_data[2278] = 33'd3933739912;
        test_addr[2279] = 50;
        test_data[2279] = 33'd2829983091;
        test_addr[2280] = 51;
        test_data[2280] = 33'd2194417863;
        test_addr[2281] = 52;
        test_data[2281] = 33'd244377089;
        test_addr[2282] = 53;
        test_data[2282] = 33'd7450953192;
        test_addr[2283] = 54;
        test_data[2283] = 33'd4032295902;
        test_addr[2284] = 55;
        test_data[2284] = 33'd7368873431;
        test_addr[2285] = 56;
        test_data[2285] = 33'd8329813561;
        test_addr[2286] = 182;
        test_data[2286] = 33'd407882722;
        test_addr[2287] = 183;
        test_data[2287] = 33'd1700753432;
        test_addr[2288] = 57;
        test_data[2288] = 33'd6467024357;
        test_addr[2289] = 58;
        test_data[2289] = 33'd3980185017;
        test_addr[2290] = 59;
        test_data[2290] = 33'd587109440;
        test_addr[2291] = 60;
        test_data[2291] = 33'd7247098673;
        test_addr[2292] = 61;
        test_data[2292] = 33'd3065752321;
        test_addr[2293] = 562;
        test_data[2293] = 33'd1942238216;
        test_addr[2294] = 563;
        test_data[2294] = 33'd3656355596;
        test_addr[2295] = 564;
        test_data[2295] = 33'd4878049514;
        test_addr[2296] = 565;
        test_data[2296] = 33'd1142270682;
        test_addr[2297] = 566;
        test_data[2297] = 33'd3267954081;
        test_addr[2298] = 567;
        test_data[2298] = 33'd6667631106;
        test_addr[2299] = 568;
        test_data[2299] = 33'd6697373523;
        test_addr[2300] = 62;
        test_data[2300] = 33'd3712003529;
        test_addr[2301] = 63;
        test_data[2301] = 33'd8219500297;
        test_addr[2302] = 64;
        test_data[2302] = 33'd3007627993;
        test_addr[2303] = 65;
        test_data[2303] = 33'd1673314307;
        test_addr[2304] = 66;
        test_data[2304] = 33'd333749771;
        test_addr[2305] = 67;
        test_data[2305] = 33'd283800910;
        test_addr[2306] = 68;
        test_data[2306] = 33'd7138449587;
        test_addr[2307] = 838;
        test_data[2307] = 33'd3624299934;
        test_addr[2308] = 839;
        test_data[2308] = 33'd2174987116;
        test_addr[2309] = 840;
        test_data[2309] = 33'd6978423349;
        test_addr[2310] = 841;
        test_data[2310] = 33'd1980186126;
        test_addr[2311] = 842;
        test_data[2311] = 33'd3536331538;
        test_addr[2312] = 843;
        test_data[2312] = 33'd1817785861;
        test_addr[2313] = 844;
        test_data[2313] = 33'd2938986312;
        test_addr[2314] = 69;
        test_data[2314] = 33'd8166525102;
        test_addr[2315] = 70;
        test_data[2315] = 33'd2063300234;
        test_addr[2316] = 71;
        test_data[2316] = 33'd5192888066;
        test_addr[2317] = 72;
        test_data[2317] = 33'd2736407674;
        test_addr[2318] = 73;
        test_data[2318] = 33'd5911311404;
        test_addr[2319] = 541;
        test_data[2319] = 33'd1842778203;
        test_addr[2320] = 542;
        test_data[2320] = 33'd3693452330;
        test_addr[2321] = 543;
        test_data[2321] = 33'd7707539472;
        test_addr[2322] = 544;
        test_data[2322] = 33'd118999468;
        test_addr[2323] = 545;
        test_data[2323] = 33'd3588739236;
        test_addr[2324] = 546;
        test_data[2324] = 33'd717909476;
        test_addr[2325] = 547;
        test_data[2325] = 33'd1656097789;
        test_addr[2326] = 548;
        test_data[2326] = 33'd3975122350;
        test_addr[2327] = 549;
        test_data[2327] = 33'd7565630825;
        test_addr[2328] = 550;
        test_data[2328] = 33'd6669382584;
        test_addr[2329] = 74;
        test_data[2329] = 33'd1226571034;
        test_addr[2330] = 75;
        test_data[2330] = 33'd1317445743;
        test_addr[2331] = 76;
        test_data[2331] = 33'd2183571412;
        test_addr[2332] = 77;
        test_data[2332] = 33'd1951277074;
        test_addr[2333] = 8;
        test_data[2333] = 33'd4074274575;
        test_addr[2334] = 9;
        test_data[2334] = 33'd5318617022;
        test_addr[2335] = 10;
        test_data[2335] = 33'd2770097472;
        test_addr[2336] = 11;
        test_data[2336] = 33'd4191856559;
        test_addr[2337] = 12;
        test_data[2337] = 33'd290304978;
        test_addr[2338] = 13;
        test_data[2338] = 33'd6860166402;
        test_addr[2339] = 78;
        test_data[2339] = 33'd3938077862;
        test_addr[2340] = 79;
        test_data[2340] = 33'd5734068344;
        test_addr[2341] = 80;
        test_data[2341] = 33'd1340395370;
        test_addr[2342] = 81;
        test_data[2342] = 33'd3320844183;
        test_addr[2343] = 699;
        test_data[2343] = 33'd2973118482;
        test_addr[2344] = 700;
        test_data[2344] = 33'd968388609;
        test_addr[2345] = 701;
        test_data[2345] = 33'd835744670;
        test_addr[2346] = 702;
        test_data[2346] = 33'd1564728561;
        test_addr[2347] = 703;
        test_data[2347] = 33'd1255659046;
        test_addr[2348] = 704;
        test_data[2348] = 33'd7128549271;
        test_addr[2349] = 705;
        test_data[2349] = 33'd1911257944;
        test_addr[2350] = 706;
        test_data[2350] = 33'd3521378079;
        test_addr[2351] = 82;
        test_data[2351] = 33'd2763428529;
        test_addr[2352] = 83;
        test_data[2352] = 33'd1828590022;
        test_addr[2353] = 84;
        test_data[2353] = 33'd1081301073;
        test_addr[2354] = 189;
        test_data[2354] = 33'd6045097381;
        test_addr[2355] = 190;
        test_data[2355] = 33'd2886127342;
        test_addr[2356] = 191;
        test_data[2356] = 33'd1659134554;
        test_addr[2357] = 85;
        test_data[2357] = 33'd725363894;
        test_addr[2358] = 345;
        test_data[2358] = 33'd209889135;
        test_addr[2359] = 346;
        test_data[2359] = 33'd6867045953;
        test_addr[2360] = 347;
        test_data[2360] = 33'd4097960042;
        test_addr[2361] = 348;
        test_data[2361] = 33'd3314453200;
        test_addr[2362] = 349;
        test_data[2362] = 33'd2590479583;
        test_addr[2363] = 350;
        test_data[2363] = 33'd1343466654;
        test_addr[2364] = 351;
        test_data[2364] = 33'd7055051613;
        test_addr[2365] = 352;
        test_data[2365] = 33'd8235940044;
        test_addr[2366] = 353;
        test_data[2366] = 33'd469648569;
        test_addr[2367] = 354;
        test_data[2367] = 33'd7916492652;
        test_addr[2368] = 355;
        test_data[2368] = 33'd7071808034;
        test_addr[2369] = 356;
        test_data[2369] = 33'd1186428617;
        test_addr[2370] = 357;
        test_data[2370] = 33'd1851805845;
        test_addr[2371] = 358;
        test_data[2371] = 33'd8522826677;
        test_addr[2372] = 359;
        test_data[2372] = 33'd7049015708;
        test_addr[2373] = 360;
        test_data[2373] = 33'd771623211;
        test_addr[2374] = 361;
        test_data[2374] = 33'd7456681815;
        test_addr[2375] = 362;
        test_data[2375] = 33'd2751591009;
        test_addr[2376] = 363;
        test_data[2376] = 33'd3362159751;
        test_addr[2377] = 86;
        test_data[2377] = 33'd6974646493;
        test_addr[2378] = 87;
        test_data[2378] = 33'd597900638;
        test_addr[2379] = 88;
        test_data[2379] = 33'd6434858146;
        test_addr[2380] = 89;
        test_data[2380] = 33'd461104171;
        test_addr[2381] = 126;
        test_data[2381] = 33'd4195730453;
        test_addr[2382] = 127;
        test_data[2382] = 33'd676159653;
        test_addr[2383] = 128;
        test_data[2383] = 33'd1760199638;
        test_addr[2384] = 129;
        test_data[2384] = 33'd652071928;
        test_addr[2385] = 130;
        test_data[2385] = 33'd4757220854;
        test_addr[2386] = 131;
        test_data[2386] = 33'd7837093478;
        test_addr[2387] = 132;
        test_data[2387] = 33'd5047035764;
        test_addr[2388] = 133;
        test_data[2388] = 33'd4531394821;
        test_addr[2389] = 90;
        test_data[2389] = 33'd43380869;
        test_addr[2390] = 914;
        test_data[2390] = 33'd6212678470;
        test_addr[2391] = 915;
        test_data[2391] = 33'd1563133648;
        test_addr[2392] = 91;
        test_data[2392] = 33'd6283394858;
        test_addr[2393] = 92;
        test_data[2393] = 33'd5838819041;
        test_addr[2394] = 93;
        test_data[2394] = 33'd7212328572;
        test_addr[2395] = 94;
        test_data[2395] = 33'd4213193887;
        test_addr[2396] = 95;
        test_data[2396] = 33'd610452162;
        test_addr[2397] = 96;
        test_data[2397] = 33'd3730512133;
        test_addr[2398] = 97;
        test_data[2398] = 33'd654962339;
        test_addr[2399] = 98;
        test_data[2399] = 33'd2789486256;
        test_addr[2400] = 99;
        test_data[2400] = 33'd1718939551;
        test_addr[2401] = 100;
        test_data[2401] = 33'd3845605637;
        test_addr[2402] = 789;
        test_data[2402] = 33'd4672343216;
        test_addr[2403] = 790;
        test_data[2403] = 33'd7749321566;
        test_addr[2404] = 791;
        test_data[2404] = 33'd206378386;
        test_addr[2405] = 792;
        test_data[2405] = 33'd4001250463;
        test_addr[2406] = 793;
        test_data[2406] = 33'd1013045164;
        test_addr[2407] = 794;
        test_data[2407] = 33'd5142231792;
        test_addr[2408] = 795;
        test_data[2408] = 33'd4412406508;
        test_addr[2409] = 796;
        test_data[2409] = 33'd3245915395;
        test_addr[2410] = 797;
        test_data[2410] = 33'd7051317930;
        test_addr[2411] = 798;
        test_data[2411] = 33'd3084085916;
        test_addr[2412] = 799;
        test_data[2412] = 33'd6320175770;
        test_addr[2413] = 800;
        test_data[2413] = 33'd4487684769;
        test_addr[2414] = 801;
        test_data[2414] = 33'd2873799072;
        test_addr[2415] = 802;
        test_data[2415] = 33'd4906220577;
        test_addr[2416] = 803;
        test_data[2416] = 33'd3660731959;
        test_addr[2417] = 804;
        test_data[2417] = 33'd3876585234;
        test_addr[2418] = 805;
        test_data[2418] = 33'd341095953;
        test_addr[2419] = 806;
        test_data[2419] = 33'd1803781852;
        test_addr[2420] = 807;
        test_data[2420] = 33'd7694975391;
        test_addr[2421] = 808;
        test_data[2421] = 33'd3811340329;
        test_addr[2422] = 809;
        test_data[2422] = 33'd2346369745;
        test_addr[2423] = 810;
        test_data[2423] = 33'd848075204;
        test_addr[2424] = 101;
        test_data[2424] = 33'd669798772;
        test_addr[2425] = 102;
        test_data[2425] = 33'd5180495055;
        test_addr[2426] = 103;
        test_data[2426] = 33'd3242132899;
        test_addr[2427] = 104;
        test_data[2427] = 33'd4408725814;
        test_addr[2428] = 105;
        test_data[2428] = 33'd4872318557;
        test_addr[2429] = 106;
        test_data[2429] = 33'd5999594103;
        test_addr[2430] = 107;
        test_data[2430] = 33'd6191521170;
        test_addr[2431] = 108;
        test_data[2431] = 33'd4486198119;
        test_addr[2432] = 109;
        test_data[2432] = 33'd6418303212;
        test_addr[2433] = 110;
        test_data[2433] = 33'd1563193765;
        test_addr[2434] = 111;
        test_data[2434] = 33'd59269632;
        test_addr[2435] = 112;
        test_data[2435] = 33'd26118987;
        test_addr[2436] = 113;
        test_data[2436] = 33'd124869335;
        test_addr[2437] = 114;
        test_data[2437] = 33'd263631887;
        test_addr[2438] = 115;
        test_data[2438] = 33'd2227853741;
        test_addr[2439] = 116;
        test_data[2439] = 33'd2133211513;
        test_addr[2440] = 117;
        test_data[2440] = 33'd8266338300;
        test_addr[2441] = 118;
        test_data[2441] = 33'd2838500611;
        test_addr[2442] = 119;
        test_data[2442] = 33'd5243636967;
        test_addr[2443] = 740;
        test_data[2443] = 33'd2567066062;
        test_addr[2444] = 741;
        test_data[2444] = 33'd2013379092;
        test_addr[2445] = 742;
        test_data[2445] = 33'd546339758;
        test_addr[2446] = 743;
        test_data[2446] = 33'd2720583043;
        test_addr[2447] = 744;
        test_data[2447] = 33'd4202166401;
        test_addr[2448] = 745;
        test_data[2448] = 33'd6791455369;
        test_addr[2449] = 746;
        test_data[2449] = 33'd6824276551;
        test_addr[2450] = 747;
        test_data[2450] = 33'd4029219969;
        test_addr[2451] = 748;
        test_data[2451] = 33'd5257252233;
        test_addr[2452] = 749;
        test_data[2452] = 33'd7392341134;
        test_addr[2453] = 120;
        test_data[2453] = 33'd8582130622;
        test_addr[2454] = 121;
        test_data[2454] = 33'd6169050649;
        test_addr[2455] = 122;
        test_data[2455] = 33'd3741684855;
        test_addr[2456] = 123;
        test_data[2456] = 33'd2458661410;
        test_addr[2457] = 124;
        test_data[2457] = 33'd2861445713;
        test_addr[2458] = 125;
        test_data[2458] = 33'd7188570028;
        test_addr[2459] = 126;
        test_data[2459] = 33'd4325905082;
        test_addr[2460] = 127;
        test_data[2460] = 33'd676159653;
        test_addr[2461] = 128;
        test_data[2461] = 33'd1760199638;
        test_addr[2462] = 129;
        test_data[2462] = 33'd652071928;
        test_addr[2463] = 185;
        test_data[2463] = 33'd845095807;
        test_addr[2464] = 186;
        test_data[2464] = 33'd621023615;
        test_addr[2465] = 187;
        test_data[2465] = 33'd6755780818;
        test_addr[2466] = 188;
        test_data[2466] = 33'd4951923185;
        test_addr[2467] = 189;
        test_data[2467] = 33'd1750130085;
        test_addr[2468] = 190;
        test_data[2468] = 33'd2886127342;
        test_addr[2469] = 191;
        test_data[2469] = 33'd1659134554;
        test_addr[2470] = 192;
        test_data[2470] = 33'd4565635275;
        test_addr[2471] = 193;
        test_data[2471] = 33'd6526375281;
        test_addr[2472] = 194;
        test_data[2472] = 33'd6698178506;
        test_addr[2473] = 195;
        test_data[2473] = 33'd6926075967;
        test_addr[2474] = 196;
        test_data[2474] = 33'd3889204301;
        test_addr[2475] = 197;
        test_data[2475] = 33'd813799808;
        test_addr[2476] = 198;
        test_data[2476] = 33'd400801465;
        test_addr[2477] = 199;
        test_data[2477] = 33'd7327254951;
        test_addr[2478] = 200;
        test_data[2478] = 33'd3223549335;
        test_addr[2479] = 201;
        test_data[2479] = 33'd4506633782;
        test_addr[2480] = 202;
        test_data[2480] = 33'd1170319904;
        test_addr[2481] = 203;
        test_data[2481] = 33'd2685333552;
        test_addr[2482] = 204;
        test_data[2482] = 33'd3227643862;
        test_addr[2483] = 205;
        test_data[2483] = 33'd5574796376;
        test_addr[2484] = 206;
        test_data[2484] = 33'd2946247101;
        test_addr[2485] = 207;
        test_data[2485] = 33'd1368502602;
        test_addr[2486] = 208;
        test_data[2486] = 33'd1843892378;
        test_addr[2487] = 209;
        test_data[2487] = 33'd798173977;
        test_addr[2488] = 130;
        test_data[2488] = 33'd462253558;
        test_addr[2489] = 131;
        test_data[2489] = 33'd8367803512;
        test_addr[2490] = 132;
        test_data[2490] = 33'd8460158215;
        test_addr[2491] = 133;
        test_data[2491] = 33'd236427525;
        test_addr[2492] = 942;
        test_data[2492] = 33'd919749232;
        test_addr[2493] = 943;
        test_data[2493] = 33'd1010987243;
        test_addr[2494] = 944;
        test_data[2494] = 33'd5802707961;
        test_addr[2495] = 945;
        test_data[2495] = 33'd158465285;
        test_addr[2496] = 946;
        test_data[2496] = 33'd4251511846;
        test_addr[2497] = 947;
        test_data[2497] = 33'd1790299456;
        test_addr[2498] = 948;
        test_data[2498] = 33'd8574615884;
        test_addr[2499] = 949;
        test_data[2499] = 33'd7830983973;
        test_addr[2500] = 950;
        test_data[2500] = 33'd7828449895;
        test_addr[2501] = 951;
        test_data[2501] = 33'd5605359386;
        test_addr[2502] = 952;
        test_data[2502] = 33'd4040559479;
        test_addr[2503] = 953;
        test_data[2503] = 33'd7164528210;
        test_addr[2504] = 954;
        test_data[2504] = 33'd5241982417;
        test_addr[2505] = 955;
        test_data[2505] = 33'd2159617400;
        test_addr[2506] = 956;
        test_data[2506] = 33'd922515263;
        test_addr[2507] = 957;
        test_data[2507] = 33'd3725935089;
        test_addr[2508] = 958;
        test_data[2508] = 33'd1131678623;
        test_addr[2509] = 134;
        test_data[2509] = 33'd2903040825;
        test_addr[2510] = 135;
        test_data[2510] = 33'd2176215843;
        test_addr[2511] = 136;
        test_data[2511] = 33'd6600150322;
        test_addr[2512] = 137;
        test_data[2512] = 33'd2464351703;
        test_addr[2513] = 138;
        test_data[2513] = 33'd6883526884;
        test_addr[2514] = 139;
        test_data[2514] = 33'd3600776137;
        test_addr[2515] = 140;
        test_data[2515] = 33'd3314446855;
        test_addr[2516] = 141;
        test_data[2516] = 33'd1108123326;
        test_addr[2517] = 142;
        test_data[2517] = 33'd4967755551;
        test_addr[2518] = 230;
        test_data[2518] = 33'd1628247242;
        test_addr[2519] = 143;
        test_data[2519] = 33'd5579527672;
        test_addr[2520] = 144;
        test_data[2520] = 33'd5760832867;
        test_addr[2521] = 145;
        test_data[2521] = 33'd1611631270;
        test_addr[2522] = 146;
        test_data[2522] = 33'd3958907471;
        test_addr[2523] = 147;
        test_data[2523] = 33'd3396137010;
        test_addr[2524] = 148;
        test_data[2524] = 33'd7833007090;
        test_addr[2525] = 149;
        test_data[2525] = 33'd6862555161;
        test_addr[2526] = 150;
        test_data[2526] = 33'd2726814038;
        test_addr[2527] = 151;
        test_data[2527] = 33'd6037232232;
        test_addr[2528] = 152;
        test_data[2528] = 33'd2716444339;
        test_addr[2529] = 153;
        test_data[2529] = 33'd8277402352;
        test_addr[2530] = 154;
        test_data[2530] = 33'd1885244835;
        test_addr[2531] = 155;
        test_data[2531] = 33'd1633875019;
        test_addr[2532] = 33;
        test_data[2532] = 33'd1455572206;
        test_addr[2533] = 34;
        test_data[2533] = 33'd3084178052;
        test_addr[2534] = 35;
        test_data[2534] = 33'd273674846;
        test_addr[2535] = 36;
        test_data[2535] = 33'd3086044954;
        test_addr[2536] = 37;
        test_data[2536] = 33'd2005231466;
        test_addr[2537] = 156;
        test_data[2537] = 33'd997076171;
        test_addr[2538] = 157;
        test_data[2538] = 33'd98365346;
        test_addr[2539] = 158;
        test_data[2539] = 33'd7067084490;
        test_addr[2540] = 159;
        test_data[2540] = 33'd875991290;
        test_addr[2541] = 160;
        test_data[2541] = 33'd2802001540;
        test_addr[2542] = 161;
        test_data[2542] = 33'd8241745651;
        test_addr[2543] = 162;
        test_data[2543] = 33'd760186910;
        test_addr[2544] = 163;
        test_data[2544] = 33'd5366697875;
        test_addr[2545] = 164;
        test_data[2545] = 33'd3847429411;
        test_addr[2546] = 165;
        test_data[2546] = 33'd2933056588;
        test_addr[2547] = 166;
        test_data[2547] = 33'd5936225092;
        test_addr[2548] = 167;
        test_data[2548] = 33'd4201079425;
        test_addr[2549] = 168;
        test_data[2549] = 33'd244697080;
        test_addr[2550] = 169;
        test_data[2550] = 33'd1473150397;
        test_addr[2551] = 170;
        test_data[2551] = 33'd1712482729;
        test_addr[2552] = 171;
        test_data[2552] = 33'd151920409;
        test_addr[2553] = 172;
        test_data[2553] = 33'd1056389529;
        test_addr[2554] = 173;
        test_data[2554] = 33'd7001689933;
        test_addr[2555] = 174;
        test_data[2555] = 33'd6075104753;
        test_addr[2556] = 175;
        test_data[2556] = 33'd8554652607;
        test_addr[2557] = 176;
        test_data[2557] = 33'd2837741477;
        test_addr[2558] = 177;
        test_data[2558] = 33'd2547298871;
        test_addr[2559] = 178;
        test_data[2559] = 33'd1390194371;
        test_addr[2560] = 455;
        test_data[2560] = 33'd1395496028;
        test_addr[2561] = 456;
        test_data[2561] = 33'd3486845368;
        test_addr[2562] = 457;
        test_data[2562] = 33'd1345025748;
        test_addr[2563] = 458;
        test_data[2563] = 33'd833450510;
        test_addr[2564] = 459;
        test_data[2564] = 33'd826235681;
        test_addr[2565] = 460;
        test_data[2565] = 33'd3390313948;
        test_addr[2566] = 461;
        test_data[2566] = 33'd1580710012;
        test_addr[2567] = 462;
        test_data[2567] = 33'd3770112161;
        test_addr[2568] = 463;
        test_data[2568] = 33'd5161921250;
        test_addr[2569] = 464;
        test_data[2569] = 33'd3147145687;
        test_addr[2570] = 465;
        test_data[2570] = 33'd8207936039;
        test_addr[2571] = 466;
        test_data[2571] = 33'd8012930075;
        test_addr[2572] = 179;
        test_data[2572] = 33'd4169806564;
        test_addr[2573] = 180;
        test_data[2573] = 33'd4690062826;
        test_addr[2574] = 181;
        test_data[2574] = 33'd485480945;
        test_addr[2575] = 182;
        test_data[2575] = 33'd5565340469;
        test_addr[2576] = 183;
        test_data[2576] = 33'd7187730361;
        test_addr[2577] = 184;
        test_data[2577] = 33'd4125218622;
        test_addr[2578] = 185;
        test_data[2578] = 33'd845095807;
        test_addr[2579] = 186;
        test_data[2579] = 33'd621023615;
        test_addr[2580] = 187;
        test_data[2580] = 33'd6675617754;
        test_addr[2581] = 188;
        test_data[2581] = 33'd656955889;
        test_addr[2582] = 189;
        test_data[2582] = 33'd1750130085;
        test_addr[2583] = 190;
        test_data[2583] = 33'd7262458732;
        test_addr[2584] = 191;
        test_data[2584] = 33'd1659134554;
        test_addr[2585] = 192;
        test_data[2585] = 33'd270667979;
        test_addr[2586] = 193;
        test_data[2586] = 33'd2231407985;
        test_addr[2587] = 194;
        test_data[2587] = 33'd2403211210;
        test_addr[2588] = 195;
        test_data[2588] = 33'd7354095134;
        test_addr[2589] = 196;
        test_data[2589] = 33'd3889204301;
        test_addr[2590] = 197;
        test_data[2590] = 33'd4749917305;
        test_addr[2591] = 198;
        test_data[2591] = 33'd7351674054;
        test_addr[2592] = 199;
        test_data[2592] = 33'd8458523207;
        test_addr[2593] = 200;
        test_data[2593] = 33'd3223549335;
        test_addr[2594] = 201;
        test_data[2594] = 33'd211666486;
        test_addr[2595] = 728;
        test_data[2595] = 33'd716320088;
        test_addr[2596] = 729;
        test_data[2596] = 33'd964607519;
        test_addr[2597] = 730;
        test_data[2597] = 33'd4429803876;
        test_addr[2598] = 731;
        test_data[2598] = 33'd1618801135;
        test_addr[2599] = 202;
        test_data[2599] = 33'd1170319904;
        test_addr[2600] = 203;
        test_data[2600] = 33'd2685333552;
        test_addr[2601] = 204;
        test_data[2601] = 33'd3227643862;
        test_addr[2602] = 205;
        test_data[2602] = 33'd1279829080;
        test_addr[2603] = 206;
        test_data[2603] = 33'd2946247101;
        test_addr[2604] = 207;
        test_data[2604] = 33'd1368502602;
        test_addr[2605] = 683;
        test_data[2605] = 33'd7639702177;
        test_addr[2606] = 684;
        test_data[2606] = 33'd1377128895;
        test_addr[2607] = 685;
        test_data[2607] = 33'd992539895;
        test_addr[2608] = 686;
        test_data[2608] = 33'd626729407;
        test_addr[2609] = 687;
        test_data[2609] = 33'd2332656559;
        test_addr[2610] = 688;
        test_data[2610] = 33'd6722461291;
        test_addr[2611] = 689;
        test_data[2611] = 33'd8377619706;
        test_addr[2612] = 690;
        test_data[2612] = 33'd1799699601;
        test_addr[2613] = 691;
        test_data[2613] = 33'd3914485233;
        test_addr[2614] = 692;
        test_data[2614] = 33'd1007332425;
        test_addr[2615] = 208;
        test_data[2615] = 33'd1843892378;
        test_addr[2616] = 209;
        test_data[2616] = 33'd798173977;
        test_addr[2617] = 422;
        test_data[2617] = 33'd962672775;
        test_addr[2618] = 423;
        test_data[2618] = 33'd3728980285;
        test_addr[2619] = 424;
        test_data[2619] = 33'd1190904379;
        test_addr[2620] = 210;
        test_data[2620] = 33'd4383751672;
        test_addr[2621] = 211;
        test_data[2621] = 33'd3948687695;
        test_addr[2622] = 212;
        test_data[2622] = 33'd3897575557;
        test_addr[2623] = 213;
        test_data[2623] = 33'd1862765609;
        test_addr[2624] = 214;
        test_data[2624] = 33'd3563881117;
        test_addr[2625] = 215;
        test_data[2625] = 33'd7233857254;
        test_addr[2626] = 216;
        test_data[2626] = 33'd8254947012;
        test_addr[2627] = 217;
        test_data[2627] = 33'd2173355106;
        test_addr[2628] = 218;
        test_data[2628] = 33'd3295815568;
        test_addr[2629] = 219;
        test_data[2629] = 33'd1970268263;
        test_addr[2630] = 472;
        test_data[2630] = 33'd3807878672;
        test_addr[2631] = 220;
        test_data[2631] = 33'd872379323;
        test_addr[2632] = 221;
        test_data[2632] = 33'd2167464279;
        test_addr[2633] = 615;
        test_data[2633] = 33'd3553517321;
        test_addr[2634] = 616;
        test_data[2634] = 33'd5549490897;
        test_addr[2635] = 617;
        test_data[2635] = 33'd6192307056;
        test_addr[2636] = 618;
        test_data[2636] = 33'd2989005313;
        test_addr[2637] = 619;
        test_data[2637] = 33'd2093912685;
        test_addr[2638] = 620;
        test_data[2638] = 33'd6372253237;
        test_addr[2639] = 621;
        test_data[2639] = 33'd2716412051;
        test_addr[2640] = 222;
        test_data[2640] = 33'd8241582102;
        test_addr[2641] = 223;
        test_data[2641] = 33'd3577816117;
        test_addr[2642] = 224;
        test_data[2642] = 33'd897321249;
        test_addr[2643] = 225;
        test_data[2643] = 33'd4582598119;
        test_addr[2644] = 226;
        test_data[2644] = 33'd2431492093;
        test_addr[2645] = 227;
        test_data[2645] = 33'd144417235;
        test_addr[2646] = 228;
        test_data[2646] = 33'd5553500674;
        test_addr[2647] = 229;
        test_data[2647] = 33'd5584807331;
        test_addr[2648] = 230;
        test_data[2648] = 33'd5357567779;
        test_addr[2649] = 231;
        test_data[2649] = 33'd4886819594;
        test_addr[2650] = 232;
        test_data[2650] = 33'd7220958569;
        test_addr[2651] = 233;
        test_data[2651] = 33'd1437501823;
        test_addr[2652] = 234;
        test_data[2652] = 33'd2569948806;
        test_addr[2653] = 235;
        test_data[2653] = 33'd3950602267;
        test_addr[2654] = 667;
        test_data[2654] = 33'd7438891679;
        test_addr[2655] = 668;
        test_data[2655] = 33'd1574161429;
        test_addr[2656] = 669;
        test_data[2656] = 33'd8403144378;
        test_addr[2657] = 670;
        test_data[2657] = 33'd5188808510;
        test_addr[2658] = 671;
        test_data[2658] = 33'd8520944537;
        test_addr[2659] = 672;
        test_data[2659] = 33'd6880465147;
        test_addr[2660] = 673;
        test_data[2660] = 33'd8579974113;
        test_addr[2661] = 674;
        test_data[2661] = 33'd2390983344;
        test_addr[2662] = 675;
        test_data[2662] = 33'd2709261325;
        test_addr[2663] = 676;
        test_data[2663] = 33'd1104785019;
        test_addr[2664] = 677;
        test_data[2664] = 33'd929867826;
        test_addr[2665] = 678;
        test_data[2665] = 33'd4735885622;
        test_addr[2666] = 679;
        test_data[2666] = 33'd3807285746;
        test_addr[2667] = 680;
        test_data[2667] = 33'd3119041072;
        test_addr[2668] = 681;
        test_data[2668] = 33'd4956454003;
        test_addr[2669] = 682;
        test_data[2669] = 33'd4880512792;
        test_addr[2670] = 683;
        test_data[2670] = 33'd3344734881;
        test_addr[2671] = 684;
        test_data[2671] = 33'd8276069193;
        test_addr[2672] = 685;
        test_data[2672] = 33'd992539895;
        test_addr[2673] = 686;
        test_data[2673] = 33'd626729407;
        test_addr[2674] = 687;
        test_data[2674] = 33'd2332656559;
        test_addr[2675] = 688;
        test_data[2675] = 33'd2427493995;
        test_addr[2676] = 689;
        test_data[2676] = 33'd4082652410;
        test_addr[2677] = 690;
        test_data[2677] = 33'd1799699601;
        test_addr[2678] = 691;
        test_data[2678] = 33'd3914485233;
        test_addr[2679] = 692;
        test_data[2679] = 33'd8446681298;
        test_addr[2680] = 693;
        test_data[2680] = 33'd1755618517;
        test_addr[2681] = 694;
        test_data[2681] = 33'd1783902209;
        test_addr[2682] = 695;
        test_data[2682] = 33'd6078257667;
        test_addr[2683] = 696;
        test_data[2683] = 33'd1053390424;
        test_addr[2684] = 697;
        test_data[2684] = 33'd6660284060;
        test_addr[2685] = 698;
        test_data[2685] = 33'd3900402421;
        test_addr[2686] = 236;
        test_data[2686] = 33'd619874774;
        test_addr[2687] = 237;
        test_data[2687] = 33'd2223698292;
        test_addr[2688] = 238;
        test_data[2688] = 33'd1309914105;
        test_addr[2689] = 974;
        test_data[2689] = 33'd3837769794;
        test_addr[2690] = 239;
        test_data[2690] = 33'd2034158352;
        test_addr[2691] = 240;
        test_data[2691] = 33'd1564295992;
        test_addr[2692] = 241;
        test_data[2692] = 33'd2634952013;
        test_addr[2693] = 242;
        test_data[2693] = 33'd8481990328;
        test_addr[2694] = 243;
        test_data[2694] = 33'd7575132489;
        test_addr[2695] = 244;
        test_data[2695] = 33'd3986444448;
        test_addr[2696] = 245;
        test_data[2696] = 33'd715123240;
        test_addr[2697] = 246;
        test_data[2697] = 33'd1555719501;
        test_addr[2698] = 247;
        test_data[2698] = 33'd4281086416;
        test_addr[2699] = 248;
        test_data[2699] = 33'd7454959941;
        test_addr[2700] = 249;
        test_data[2700] = 33'd1002837958;
        test_addr[2701] = 250;
        test_data[2701] = 33'd6129123424;
        test_addr[2702] = 251;
        test_data[2702] = 33'd1827628710;
        test_addr[2703] = 252;
        test_data[2703] = 33'd4594872903;
        test_addr[2704] = 253;
        test_data[2704] = 33'd1046892784;
        test_addr[2705] = 254;
        test_data[2705] = 33'd893686890;
        test_addr[2706] = 232;
        test_data[2706] = 33'd7843049687;
        test_addr[2707] = 233;
        test_data[2707] = 33'd7719663637;
        test_addr[2708] = 234;
        test_data[2708] = 33'd5311621639;
        test_addr[2709] = 235;
        test_data[2709] = 33'd3950602267;
        test_addr[2710] = 236;
        test_data[2710] = 33'd6481125572;
        test_addr[2711] = 237;
        test_data[2711] = 33'd2223698292;
        test_addr[2712] = 238;
        test_data[2712] = 33'd1309914105;
        test_addr[2713] = 239;
        test_data[2713] = 33'd2034158352;
        test_addr[2714] = 240;
        test_data[2714] = 33'd1564295992;
        test_addr[2715] = 241;
        test_data[2715] = 33'd7195939355;
        test_addr[2716] = 255;
        test_data[2716] = 33'd738701221;
        test_addr[2717] = 256;
        test_data[2717] = 33'd1838035664;
        test_addr[2718] = 809;
        test_data[2718] = 33'd2346369745;
        test_addr[2719] = 810;
        test_data[2719] = 33'd848075204;
        test_addr[2720] = 811;
        test_data[2720] = 33'd8052888083;
        test_addr[2721] = 812;
        test_data[2721] = 33'd3736148023;
        test_addr[2722] = 813;
        test_data[2722] = 33'd2586361486;
        test_addr[2723] = 814;
        test_data[2723] = 33'd8478724469;
        test_addr[2724] = 815;
        test_data[2724] = 33'd3769770053;
        test_addr[2725] = 816;
        test_data[2725] = 33'd7833951193;
        test_addr[2726] = 817;
        test_data[2726] = 33'd788918906;
        test_addr[2727] = 818;
        test_data[2727] = 33'd3877886931;
        test_addr[2728] = 257;
        test_data[2728] = 33'd3066856557;
        test_addr[2729] = 258;
        test_data[2729] = 33'd968192007;
        test_addr[2730] = 259;
        test_data[2730] = 33'd2066806968;
        test_addr[2731] = 260;
        test_data[2731] = 33'd3784376997;
        test_addr[2732] = 261;
        test_data[2732] = 33'd1628122850;
        test_addr[2733] = 262;
        test_data[2733] = 33'd4745303276;
        test_addr[2734] = 263;
        test_data[2734] = 33'd1168259603;
        test_addr[2735] = 264;
        test_data[2735] = 33'd8465577673;
        test_addr[2736] = 542;
        test_data[2736] = 33'd3693452330;
        test_addr[2737] = 543;
        test_data[2737] = 33'd6804060479;
        test_addr[2738] = 544;
        test_data[2738] = 33'd118999468;
        test_addr[2739] = 545;
        test_data[2739] = 33'd3588739236;
        test_addr[2740] = 546;
        test_data[2740] = 33'd717909476;
        test_addr[2741] = 547;
        test_data[2741] = 33'd1656097789;
        test_addr[2742] = 548;
        test_data[2742] = 33'd6547950255;
        test_addr[2743] = 549;
        test_data[2743] = 33'd3270663529;
        test_addr[2744] = 550;
        test_data[2744] = 33'd5383780111;
        test_addr[2745] = 551;
        test_data[2745] = 33'd3550124624;
        test_addr[2746] = 552;
        test_data[2746] = 33'd5520612073;
        test_addr[2747] = 553;
        test_data[2747] = 33'd1687299562;
        test_addr[2748] = 554;
        test_data[2748] = 33'd7354095386;
        test_addr[2749] = 555;
        test_data[2749] = 33'd7448347873;
        test_addr[2750] = 556;
        test_data[2750] = 33'd2939472687;
        test_addr[2751] = 557;
        test_data[2751] = 33'd985122537;
        test_addr[2752] = 558;
        test_data[2752] = 33'd911700634;
        test_addr[2753] = 559;
        test_data[2753] = 33'd5172396568;
        test_addr[2754] = 560;
        test_data[2754] = 33'd7300820584;
        test_addr[2755] = 561;
        test_data[2755] = 33'd5213281932;
        test_addr[2756] = 265;
        test_data[2756] = 33'd4232753553;
        test_addr[2757] = 266;
        test_data[2757] = 33'd1763155380;
        test_addr[2758] = 267;
        test_data[2758] = 33'd2666779884;
        test_addr[2759] = 268;
        test_data[2759] = 33'd878985346;
        test_addr[2760] = 269;
        test_data[2760] = 33'd3738711814;
        test_addr[2761] = 270;
        test_data[2761] = 33'd5407319706;
        test_addr[2762] = 271;
        test_data[2762] = 33'd6179324732;
        test_addr[2763] = 272;
        test_data[2763] = 33'd3903591382;
        test_addr[2764] = 273;
        test_data[2764] = 33'd2852287615;
        test_addr[2765] = 274;
        test_data[2765] = 33'd3297475855;
        test_addr[2766] = 275;
        test_data[2766] = 33'd1702449685;
        test_addr[2767] = 276;
        test_data[2767] = 33'd151084863;
        test_addr[2768] = 277;
        test_data[2768] = 33'd1313409944;
        test_addr[2769] = 278;
        test_data[2769] = 33'd7535823356;
        test_addr[2770] = 279;
        test_data[2770] = 33'd7314086138;
        test_addr[2771] = 280;
        test_data[2771] = 33'd4533129346;
        test_addr[2772] = 281;
        test_data[2772] = 33'd5882289519;
        test_addr[2773] = 282;
        test_data[2773] = 33'd7254028917;
        test_addr[2774] = 283;
        test_data[2774] = 33'd597342362;
        test_addr[2775] = 284;
        test_data[2775] = 33'd3042846807;
        test_addr[2776] = 285;
        test_data[2776] = 33'd7301526529;
        test_addr[2777] = 286;
        test_data[2777] = 33'd2730571741;
        test_addr[2778] = 287;
        test_data[2778] = 33'd4230987602;
        test_addr[2779] = 288;
        test_data[2779] = 33'd3200330683;
        test_addr[2780] = 289;
        test_data[2780] = 33'd2070000467;
        test_addr[2781] = 290;
        test_data[2781] = 33'd2990572821;
        test_addr[2782] = 257;
        test_data[2782] = 33'd3066856557;
        test_addr[2783] = 258;
        test_data[2783] = 33'd968192007;
        test_addr[2784] = 291;
        test_data[2784] = 33'd669926597;
        test_addr[2785] = 292;
        test_data[2785] = 33'd1963688468;
        test_addr[2786] = 293;
        test_data[2786] = 33'd4088931545;
        test_addr[2787] = 294;
        test_data[2787] = 33'd3937214664;
        test_addr[2788] = 295;
        test_data[2788] = 33'd4674692420;
        test_addr[2789] = 296;
        test_data[2789] = 33'd124823375;
        test_addr[2790] = 297;
        test_data[2790] = 33'd4656986776;
        test_addr[2791] = 298;
        test_data[2791] = 33'd2992906690;
        test_addr[2792] = 299;
        test_data[2792] = 33'd3630541901;
        test_addr[2793] = 300;
        test_data[2793] = 33'd1786211448;
        test_addr[2794] = 301;
        test_data[2794] = 33'd178124090;
        test_addr[2795] = 302;
        test_data[2795] = 33'd8589374918;
        test_addr[2796] = 303;
        test_data[2796] = 33'd7784190614;
        test_addr[2797] = 304;
        test_data[2797] = 33'd3927615128;
        test_addr[2798] = 305;
        test_data[2798] = 33'd1996090555;
        test_addr[2799] = 306;
        test_data[2799] = 33'd4071353466;
        test_addr[2800] = 307;
        test_data[2800] = 33'd4030103948;
        test_addr[2801] = 308;
        test_data[2801] = 33'd4922453240;
        test_addr[2802] = 309;
        test_data[2802] = 33'd1328657515;
        test_addr[2803] = 553;
        test_data[2803] = 33'd1687299562;
        test_addr[2804] = 554;
        test_data[2804] = 33'd3059128090;
        test_addr[2805] = 310;
        test_data[2805] = 33'd7219780933;
        test_addr[2806] = 311;
        test_data[2806] = 33'd3422864683;
        test_addr[2807] = 312;
        test_data[2807] = 33'd2136184510;
        test_addr[2808] = 313;
        test_data[2808] = 33'd3975800125;
        test_addr[2809] = 314;
        test_data[2809] = 33'd1771827745;
        test_addr[2810] = 315;
        test_data[2810] = 33'd1032608502;
        test_addr[2811] = 316;
        test_data[2811] = 33'd2961835101;
        test_addr[2812] = 317;
        test_data[2812] = 33'd613544344;
        test_addr[2813] = 318;
        test_data[2813] = 33'd1370421073;
        test_addr[2814] = 319;
        test_data[2814] = 33'd180363106;
        test_addr[2815] = 921;
        test_data[2815] = 33'd1245013432;
        test_addr[2816] = 922;
        test_data[2816] = 33'd7240868723;
        test_addr[2817] = 923;
        test_data[2817] = 33'd3103545132;
        test_addr[2818] = 924;
        test_data[2818] = 33'd1593791081;
        test_addr[2819] = 925;
        test_data[2819] = 33'd1313195782;
        test_addr[2820] = 926;
        test_data[2820] = 33'd347576106;
        test_addr[2821] = 927;
        test_data[2821] = 33'd4267639243;
        test_addr[2822] = 928;
        test_data[2822] = 33'd1094388041;
        test_addr[2823] = 929;
        test_data[2823] = 33'd1467497009;
        test_addr[2824] = 930;
        test_data[2824] = 33'd6414004925;
        test_addr[2825] = 931;
        test_data[2825] = 33'd1776715744;
        test_addr[2826] = 932;
        test_data[2826] = 33'd360085129;
        test_addr[2827] = 933;
        test_data[2827] = 33'd6667343922;
        test_addr[2828] = 934;
        test_data[2828] = 33'd392045396;
        test_addr[2829] = 935;
        test_data[2829] = 33'd2632191667;
        test_addr[2830] = 936;
        test_data[2830] = 33'd3408512394;
        test_addr[2831] = 937;
        test_data[2831] = 33'd6380541598;
        test_addr[2832] = 938;
        test_data[2832] = 33'd408550941;
        test_addr[2833] = 939;
        test_data[2833] = 33'd1167784344;
        test_addr[2834] = 940;
        test_data[2834] = 33'd5461679573;
        test_addr[2835] = 941;
        test_data[2835] = 33'd5057150948;
        test_addr[2836] = 942;
        test_data[2836] = 33'd919749232;
        test_addr[2837] = 943;
        test_data[2837] = 33'd1010987243;
        test_addr[2838] = 944;
        test_data[2838] = 33'd1507740665;
        test_addr[2839] = 945;
        test_data[2839] = 33'd158465285;
        test_addr[2840] = 946;
        test_data[2840] = 33'd4251511846;
        test_addr[2841] = 947;
        test_data[2841] = 33'd1790299456;
        test_addr[2842] = 948;
        test_data[2842] = 33'd4279648588;
        test_addr[2843] = 949;
        test_data[2843] = 33'd3536016677;
        test_addr[2844] = 950;
        test_data[2844] = 33'd3533482599;
        test_addr[2845] = 320;
        test_data[2845] = 33'd4010594226;
        test_addr[2846] = 321;
        test_data[2846] = 33'd4506111488;
        test_addr[2847] = 322;
        test_data[2847] = 33'd2250922743;
        test_addr[2848] = 323;
        test_data[2848] = 33'd6326753176;
        test_addr[2849] = 324;
        test_data[2849] = 33'd4124680673;
        test_addr[2850] = 623;
        test_data[2850] = 33'd4602239611;
        test_addr[2851] = 624;
        test_data[2851] = 33'd50566768;
        test_addr[2852] = 625;
        test_data[2852] = 33'd4595332734;
        test_addr[2853] = 626;
        test_data[2853] = 33'd489015939;
        test_addr[2854] = 627;
        test_data[2854] = 33'd157889119;
        test_addr[2855] = 628;
        test_data[2855] = 33'd2298215631;
        test_addr[2856] = 629;
        test_data[2856] = 33'd6779549984;
        test_addr[2857] = 630;
        test_data[2857] = 33'd129078420;
        test_addr[2858] = 631;
        test_data[2858] = 33'd5146463087;
        test_addr[2859] = 632;
        test_data[2859] = 33'd1956628422;
        test_addr[2860] = 633;
        test_data[2860] = 33'd5447732667;
        test_addr[2861] = 634;
        test_data[2861] = 33'd2429702712;
        test_addr[2862] = 635;
        test_data[2862] = 33'd1607332002;
        test_addr[2863] = 636;
        test_data[2863] = 33'd2340019269;
        test_addr[2864] = 637;
        test_data[2864] = 33'd1005752581;
        test_addr[2865] = 638;
        test_data[2865] = 33'd4136659456;
        test_addr[2866] = 639;
        test_data[2866] = 33'd86901798;
        test_addr[2867] = 325;
        test_data[2867] = 33'd7862708571;
        test_addr[2868] = 326;
        test_data[2868] = 33'd3211040190;
        test_addr[2869] = 327;
        test_data[2869] = 33'd4021375997;
        test_addr[2870] = 328;
        test_data[2870] = 33'd6489802474;
        test_addr[2871] = 720;
        test_data[2871] = 33'd7755793717;
        test_addr[2872] = 721;
        test_data[2872] = 33'd662721243;
        test_addr[2873] = 722;
        test_data[2873] = 33'd7805459547;
        test_addr[2874] = 723;
        test_data[2874] = 33'd2035228107;
        test_addr[2875] = 724;
        test_data[2875] = 33'd3488346519;
        test_addr[2876] = 725;
        test_data[2876] = 33'd4023969800;
        test_addr[2877] = 726;
        test_data[2877] = 33'd7845115935;
        test_addr[2878] = 727;
        test_data[2878] = 33'd7351930625;
        test_addr[2879] = 728;
        test_data[2879] = 33'd716320088;
        test_addr[2880] = 729;
        test_data[2880] = 33'd964607519;
        test_addr[2881] = 329;
        test_data[2881] = 33'd508970632;
        test_addr[2882] = 330;
        test_data[2882] = 33'd2871069657;
        test_addr[2883] = 331;
        test_data[2883] = 33'd3021584846;
        test_addr[2884] = 332;
        test_data[2884] = 33'd3802541065;
        test_addr[2885] = 333;
        test_data[2885] = 33'd3777587601;
        test_addr[2886] = 334;
        test_data[2886] = 33'd5686364335;
        test_addr[2887] = 335;
        test_data[2887] = 33'd3132902255;
        test_addr[2888] = 336;
        test_data[2888] = 33'd535597245;
        test_addr[2889] = 337;
        test_data[2889] = 33'd2803068549;
        test_addr[2890] = 338;
        test_data[2890] = 33'd1957293410;
        test_addr[2891] = 339;
        test_data[2891] = 33'd4595659399;
        test_addr[2892] = 523;
        test_data[2892] = 33'd1659053730;
        test_addr[2893] = 524;
        test_data[2893] = 33'd2535488802;
        test_addr[2894] = 525;
        test_data[2894] = 33'd2367555368;
        test_addr[2895] = 526;
        test_data[2895] = 33'd2518142267;
        test_addr[2896] = 527;
        test_data[2896] = 33'd5338216397;
        test_addr[2897] = 528;
        test_data[2897] = 33'd7466321197;
        test_addr[2898] = 529;
        test_data[2898] = 33'd6447168953;
        test_addr[2899] = 530;
        test_data[2899] = 33'd1192716121;
        test_addr[2900] = 531;
        test_data[2900] = 33'd591809078;
        test_addr[2901] = 532;
        test_data[2901] = 33'd4946991630;
        test_addr[2902] = 340;
        test_data[2902] = 33'd8282622553;
        test_addr[2903] = 341;
        test_data[2903] = 33'd3105826626;
        test_addr[2904] = 960;
        test_data[2904] = 33'd813414639;
        test_addr[2905] = 961;
        test_data[2905] = 33'd4498366049;
        test_addr[2906] = 962;
        test_data[2906] = 33'd3660914740;
        test_addr[2907] = 342;
        test_data[2907] = 33'd6346496058;
        test_addr[2908] = 343;
        test_data[2908] = 33'd3938949624;
        test_addr[2909] = 344;
        test_data[2909] = 33'd3293331081;
        test_addr[2910] = 345;
        test_data[2910] = 33'd5819449830;
        test_addr[2911] = 346;
        test_data[2911] = 33'd2572078657;
        test_addr[2912] = 347;
        test_data[2912] = 33'd4097960042;
        test_addr[2913] = 348;
        test_data[2913] = 33'd7524987529;
        test_addr[2914] = 349;
        test_data[2914] = 33'd2590479583;
        test_addr[2915] = 350;
        test_data[2915] = 33'd1343466654;
        test_addr[2916] = 613;
        test_data[2916] = 33'd3917815039;
        test_addr[2917] = 351;
        test_data[2917] = 33'd2760084317;
        test_addr[2918] = 352;
        test_data[2918] = 33'd3940972748;
        test_addr[2919] = 353;
        test_data[2919] = 33'd5217438905;
        test_addr[2920] = 354;
        test_data[2920] = 33'd4787764898;
        test_addr[2921] = 355;
        test_data[2921] = 33'd2776840738;
        test_addr[2922] = 356;
        test_data[2922] = 33'd1186428617;
        test_addr[2923] = 357;
        test_data[2923] = 33'd1851805845;
        test_addr[2924] = 358;
        test_data[2924] = 33'd4227859381;
        test_addr[2925] = 359;
        test_data[2925] = 33'd5920327461;
        test_addr[2926] = 360;
        test_data[2926] = 33'd771623211;
        test_addr[2927] = 361;
        test_data[2927] = 33'd7730528321;
        test_addr[2928] = 362;
        test_data[2928] = 33'd2751591009;
        test_addr[2929] = 363;
        test_data[2929] = 33'd3362159751;
        test_addr[2930] = 364;
        test_data[2930] = 33'd4091092656;
        test_addr[2931] = 365;
        test_data[2931] = 33'd3157196662;
        test_addr[2932] = 366;
        test_data[2932] = 33'd2904869292;
        test_addr[2933] = 367;
        test_data[2933] = 33'd7350813094;
        test_addr[2934] = 368;
        test_data[2934] = 33'd1594529834;
        test_addr[2935] = 369;
        test_data[2935] = 33'd1912926533;
        test_addr[2936] = 370;
        test_data[2936] = 33'd4639411115;
        test_addr[2937] = 371;
        test_data[2937] = 33'd1096870004;
        test_addr[2938] = 372;
        test_data[2938] = 33'd1927727626;
        test_addr[2939] = 373;
        test_data[2939] = 33'd3498474298;
        test_addr[2940] = 374;
        test_data[2940] = 33'd149363693;
        test_addr[2941] = 375;
        test_data[2941] = 33'd7014182649;
        test_addr[2942] = 376;
        test_data[2942] = 33'd736569085;
        test_addr[2943] = 377;
        test_data[2943] = 33'd4792875971;
        test_addr[2944] = 378;
        test_data[2944] = 33'd506127913;
        test_addr[2945] = 379;
        test_data[2945] = 33'd8199296524;
        test_addr[2946] = 380;
        test_data[2946] = 33'd2614266083;
        test_addr[2947] = 381;
        test_data[2947] = 33'd5613258948;
        test_addr[2948] = 382;
        test_data[2948] = 33'd2994681403;
        test_addr[2949] = 383;
        test_data[2949] = 33'd461073433;
        test_addr[2950] = 384;
        test_data[2950] = 33'd739005625;
        test_addr[2951] = 495;
        test_data[2951] = 33'd759490144;
        test_addr[2952] = 496;
        test_data[2952] = 33'd667303173;
        test_addr[2953] = 497;
        test_data[2953] = 33'd6244579413;
        test_addr[2954] = 385;
        test_data[2954] = 33'd698224158;
        test_addr[2955] = 386;
        test_data[2955] = 33'd6848058184;
        test_addr[2956] = 931;
        test_data[2956] = 33'd7962799624;
        test_addr[2957] = 932;
        test_data[2957] = 33'd360085129;
        test_addr[2958] = 933;
        test_data[2958] = 33'd7527200989;
        test_addr[2959] = 934;
        test_data[2959] = 33'd392045396;
        test_addr[2960] = 935;
        test_data[2960] = 33'd5032966871;
        test_addr[2961] = 387;
        test_data[2961] = 33'd140765230;
        test_addr[2962] = 388;
        test_data[2962] = 33'd4211620500;
        test_addr[2963] = 389;
        test_data[2963] = 33'd1130499402;
        test_addr[2964] = 390;
        test_data[2964] = 33'd2928158067;
        test_addr[2965] = 391;
        test_data[2965] = 33'd4972572383;
        test_addr[2966] = 392;
        test_data[2966] = 33'd10599762;
        test_addr[2967] = 243;
        test_data[2967] = 33'd3280165193;
        test_addr[2968] = 244;
        test_data[2968] = 33'd3986444448;
        test_addr[2969] = 245;
        test_data[2969] = 33'd7330720011;
        test_addr[2970] = 246;
        test_data[2970] = 33'd1555719501;
        test_addr[2971] = 247;
        test_data[2971] = 33'd8151785655;
        test_addr[2972] = 248;
        test_data[2972] = 33'd3159992645;
        test_addr[2973] = 249;
        test_data[2973] = 33'd1002837958;
        test_addr[2974] = 250;
        test_data[2974] = 33'd7450795206;
        test_addr[2975] = 251;
        test_data[2975] = 33'd1827628710;
        test_addr[2976] = 252;
        test_data[2976] = 33'd299905607;
        test_addr[2977] = 393;
        test_data[2977] = 33'd1215078312;
        test_addr[2978] = 394;
        test_data[2978] = 33'd3640178936;
        test_addr[2979] = 395;
        test_data[2979] = 33'd4037953191;
        test_addr[2980] = 396;
        test_data[2980] = 33'd7437192972;
        test_addr[2981] = 397;
        test_data[2981] = 33'd8119819531;
        test_addr[2982] = 398;
        test_data[2982] = 33'd7618506640;
        test_addr[2983] = 399;
        test_data[2983] = 33'd798523023;
        test_addr[2984] = 400;
        test_data[2984] = 33'd12061985;
        test_addr[2985] = 544;
        test_data[2985] = 33'd6517969974;
        test_addr[2986] = 545;
        test_data[2986] = 33'd3588739236;
        test_addr[2987] = 546;
        test_data[2987] = 33'd4926311107;
        test_addr[2988] = 401;
        test_data[2988] = 33'd1367308988;
        test_addr[2989] = 402;
        test_data[2989] = 33'd3328109157;
        test_addr[2990] = 403;
        test_data[2990] = 33'd1931821484;
        test_addr[2991] = 404;
        test_data[2991] = 33'd1720976526;
        test_addr[2992] = 1020;
        test_data[2992] = 33'd1661472402;
        test_addr[2993] = 1021;
        test_data[2993] = 33'd229156893;
        test_addr[2994] = 1022;
        test_data[2994] = 33'd657762763;
        test_addr[2995] = 1023;
        test_data[2995] = 33'd2095860060;
        test_addr[2996] = 0;
        test_data[2996] = 33'd597582581;
        test_addr[2997] = 1;
        test_data[2997] = 33'd365228161;
        test_addr[2998] = 2;
        test_data[2998] = 33'd244488320;
        test_addr[2999] = 3;
        test_data[2999] = 33'd2009627834;

    end
endmodule
